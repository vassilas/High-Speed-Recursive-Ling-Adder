// Stage 1
//--------------------------------------------------------------------------------------
module J64_stage_1(a, b, g, p, x, R1, Q1);
//
//
//
    input [63:0]a ;
    input [63:0]b ;
    output [63:0]g ;
    output [63:0]p ;
    output [63:0]x ;
    output [63:0]R1 ;
    output [63:0]Q1 ;
    
    
    assign p[63:0] = a[63:0] | b[63:0] ;
    assign g[63:0] = a[63:0] & b[63:0] ;
    assign x[63:0] = a[63:0] ^ b[63:0] ;   

    
    assign R1[63:0] = g[63:0] | {g[62:0],g[63]};
    assign Q1[63:0] = p[63:0] & {p[62:0],p[63]} ;
    
endmodule


// Stage 2
//--------------------------------------------------------------------------------------
module J64_stage_2(R1, Q1, R2, Q2);
//
//
//
    input [63:0]R1;
    input [63:0]Q1;
    output [63:0]R2;
    output [63:0]Q2;

    assign R2[63:0] = R1[63:0] | {R1[61:0],R1[63:62]} | {Q1[60:0],Q1[63:61]} & {R1[59:0],R1[63:60]} | {Q1[60:0],Q1[63:61]}&{Q1[58:0],Q1[63:59]}&{R1[57:0],R1[63:58]} ;
    assign Q2[63:0] = Q1[63:0] & {Q1[61:0],Q1[63:62]} & {Q1[59:0],Q1[63:60]} & ({R1[58:0],R1[63:59]} | {Q1[57:0],Q1[63:58]});

    
endmodule



// Stage 3
//--------------------------------------------------------------------------------------
module J64_stage_3(R2, Q2, R3, Q3);
//
//
//
    input [63:0]R2;
    input [63:0]Q2;
    output [63:0]R3;
    output [63:0]Q3;

    assign R3[63:0] = R2[63:0] | {R2[55:0],R2[63:56]} | {Q2[52:0],Q2[63:53]} & {R2[47:0],R2[63:48]} | {Q2[52:0],Q2[63:53]} & {Q2[44:0],Q2[63:45]} & {R2[39:0],R2[63:40]} ;
    assign Q3[63:0] = Q2[63:0] & {Q2[55:0],Q2[63:56]} & {Q2[47:0],Q2[63:48]} & ( {R2[42:0],R2[63:43]}  |  {Q2[39:0],Q2[63:40]} ) ;
    
endmodule



// Stage 4
//--------------------------------------------------------------------------------------
module J64_stage_4(R3, Q3, R4);
//
//
//
    input [63:0]R3;
    input [63:0]Q3;
    output [63:0]R4;

    assign R4[63:0] = R3[63:0] | ( {Q3[52:0],Q3[63:53]} & {R3[31:0],R3[63:32]} ) ;
    
endmodule


// D recursion
//--------------------------------------------------------------------------------------
module J64_D_recursion(p,g,x,R2,Q2,D,xD);
    input [63:0]p;
    input [63:0]g;
    input [63:0]x;
    input [63:0]Q2;
    input [63:0]R2;
    output [63:0]D;
    output [63:0]xD;    
    
    wire [63:0]D_r;
    
    assign D_r[63:0] = g[63:0] | p[63:0]&{g[62:0],g[63]} | p[63:0]&{p[62:0],p[63]}&{p[61:0],p[63:62]} ;
    
    assign D[63:0] = D_r[63:0] & ( R2[63:0] | {Q2[60:0],Q2[63:61]} ) ;
    assign xD[63:0] = x[63:0] ^ {D[62:0],D[63]} ;
endmodule


// Adder
//--------------------------------------------------------------------------------------
module J64_adder(a, b, sum);
//
//
//
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    
    wire [63:0] g ;
    wire [63:0] p ;
    wire [63:0] x ;    
    wire [63:0] R1 ;
    wire [63:0] R2 ;
    wire [63:0] R3 ;
    wire [63:0] R4 ;
    wire [63:0] Q1 ;
    wire [63:0] Q2 ;
    wire [63:0] Q3 ;
    wire [63:0] D ;
    wire [63:0] xD ;
    
    J64_stage_1 CUT1(a, b, g, p, x, R1, Q1);
    J64_stage_2 CUT2(R1, Q1, R2, Q2);
    J64_stage_3 CUT3(R2,Q2,R3,Q3);
    J64_stage_4 CUT4(R3, Q3, R4);
    J64_D_recursion CUT5(p,g,x,R2,Q2,D,xD);
    
    assign sum[63:0] = ~{R4[62:0],R4[63]} & x[63:0] | {R4[62:0],R4[63]} & xD[63:0] ;

    
endmodule










// Architecture 4x4x4
//--------------------------------------------------------------------------------------

// Stage 1
//--------------------------------------------------------------------------------------
module J4x4x4_stage_1(a, b, g, p, x, R1, Q1, D1);
//
//
//
    input [63:0]a ;
    input [63:0]b ;
    output [63:0]g ;
    output [63:0]p ;
    output [63:0]x ;
    output [63:0]R1 ;
    output [63:0]Q1 ;
    output [63:0]D1 ;    
    
    assign p[63:0] = a[63:0] | b[63:0] ;
    assign g[63:0] = a[63:0] & b[63:0] ;
    assign x[63:0] = a[63:0] ^ b[63:0] ;   

    
    assign R1[63:0] =   g[63:0] | 
                        {g[62:0],g[63]} | 
                        {p[62:0],p[63]} & {g[61:0],g[63:62]} | 
                        {p[62:0],p[63]} & {p[61:0],p[63:62]} & {g[60:0],g[63:61]} ;
                        
                        
    assign Q1[63:0] =   p[63:0] & 
                        {p[62:0],p[63]} & 
                        {p[61:0],p[63:62]} & 
                        {p[60:0],p[63:61]}  ;

    assign D1[63:0] = p[63:0] & (   g[63:0] | 
                                    {g[62:0],g[63]} |  
                                    {p[62:0],p[63]} & {g[61:0],g[63:62]} | 
                                    {p[62:0],p[63]} & {p[61:0],p[63:62]} 
                                ) ;
                        
endmodule


// Stage 2
//--------------------------------------------------------------------------------------
module J4x4x4_stage_2(R1, Q1, D1, R2, Q2, D2);
//
//
//
    input [63:0]R1 ;
    input [63:0]Q1 ;
    input [63:0]D1 ;
    output [63:0]R2 ;
    output [63:0]Q2 ;
    output [63:0]D2 ;    
  

    
    assign R2[63:0] =   R1[63:0] |
                        {R1[59:0],R1[63:60]} |
                        {Q1[58:0],Q1[63:59]} & {R1[55:0],R1[63:56]} |
                        {Q1[58:0],Q1[63:59]} & {Q1[54:0],Q1[63:55]} & {R1[51:0],R1[63:52]} ;
    
    assign Q2[63:0] =  Q1[63:0] & {Q1[59:0],Q1[63:60]} & {Q1[55:0],Q1[63:56]} & ( {R1[52:0],R1[63:53]} | {Q1[51:0],Q1[63:52]}  ) ;
    
    assign D2[63:0] = D1[63:0] & (  R1[63:0] | {Q1[62:0],Q1[63]} ) ;
endmodule


// Stage 3
//--------------------------------------------------------------------------------------
module J4x4x4_stage_3(R2, Q2, x, D2, R3, xD);
//
//
//
    input [63:0]R2 ;
    input [63:0]Q2 ;
    input [63:0]x ;      
    input [63:0]D2 ;
    output [63:0]R3 ;
    output [63:0]xD ;
    
    wire [63:0]D ;
    
    assign R3[63:0] =   R2[63:0] |
                        {R2[47:0],R2[63:48]} |
                        {Q2[42:0],Q2[63:43]} & {R2[31:0],R2[63:32]} |
                        {Q2[42:0],Q2[63:43]} & {Q2[26:0],Q2[63:27]} & {R2[15:0],R2[63:16]} ;

    assign D[63:0] = D2[63:0] & (  R2[63:0] |  {Q2[58:0],Q2[63:59]} ) ;
    
    assign xD[63:0] = x[63:0] ^ {D[62:0],D[63]} ; 
    
endmodule






// Adder 4x4x4
//--------------------------------------------------------------------------------------
module J4x4x4_adder(a, b, sum);
//
//
//
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    

    wire [63:0] p ; 
    wire [63:0] g ;     
    wire [63:0] x ;    
    wire [63:0] R1 ;
    wire [63:0] R2 ;
    wire [63:0] R3 ;
    wire [63:0] Q1 ;
    wire [63:0] Q2 ;
    wire [63:0] D1 ;
    wire [63:0] D2 ;
    wire [63:0] xD ;
    
    J4x4x4_stage_1 CUT1(a, b, g, p, x, R1, Q1, D1);
    J4x4x4_stage_2 CUT2(R1, Q1, D1, R2, Q2, D2);
    J4x4x4_stage_3 CUT3(R2, Q2, x, D2, R3, xD);
    
    
    
    
    assign sum[63:0] = ~{R3[62:0],R3[63]} & x[63:0] | {R3[62:0],R3[63]} & xD[63:0] ;

    
endmodule


