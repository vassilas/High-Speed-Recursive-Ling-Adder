module L64_node_adder(a, b, sum);
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    wire [63:0]g ;
    wire [63:0]p ;
    wire [63:0]x ;
    wire [63:0]H1 ;
    wire [63:0]H2 ;
    wire [63:0]H3 ;
    wire [63:0]Pr1 ;
    wire [63:0]Pr2 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;
    _gpx _gpx_16	(a[16],	b[16],	g[16], 	p[16], 	x[16]) ;
    _gpx _gpx_17	(a[17],	b[17],	g[17], 	p[17], 	x[17]) ;
    _gpx _gpx_18	(a[18],	b[18],	g[18], 	p[18], 	x[18]) ;
    _gpx _gpx_19	(a[19],	b[19],	g[19], 	p[19], 	x[19]) ;
    _gpx _gpx_20	(a[20],	b[20],	g[20], 	p[20], 	x[20]) ;
    _gpx _gpx_21	(a[21],	b[21],	g[21], 	p[21], 	x[21]) ;
    _gpx _gpx_22	(a[22],	b[22],	g[22], 	p[22], 	x[22]) ;
    _gpx _gpx_23	(a[23],	b[23],	g[23], 	p[23], 	x[23]) ;
    _gpx _gpx_24	(a[24],	b[24],	g[24], 	p[24], 	x[24]) ;
    _gpx _gpx_25	(a[25],	b[25],	g[25], 	p[25], 	x[25]) ;
    _gpx _gpx_26	(a[26],	b[26],	g[26], 	p[26], 	x[26]) ;
    _gpx _gpx_27	(a[27],	b[27],	g[27], 	p[27], 	x[27]) ;
    _gpx _gpx_28	(a[28],	b[28],	g[28], 	p[28], 	x[28]) ;
    _gpx _gpx_29	(a[29],	b[29],	g[29], 	p[29], 	x[29]) ;
    _gpx _gpx_30	(a[30],	b[30],	g[30], 	p[30], 	x[30]) ;
    _gpx _gpx_31	(a[31],	b[31],	g[31], 	p[31], 	x[31]) ;
    _gpx _gpx_32	(a[32],	b[32],	g[32], 	p[32], 	x[32]) ;
    _gpx _gpx_33	(a[33],	b[33],	g[33], 	p[33], 	x[33]) ;
    _gpx _gpx_34	(a[34],	b[34],	g[34], 	p[34], 	x[34]) ;
    _gpx _gpx_35	(a[35],	b[35],	g[35], 	p[35], 	x[35]) ;
    _gpx _gpx_36	(a[36],	b[36],	g[36], 	p[36], 	x[36]) ;
    _gpx _gpx_37	(a[37],	b[37],	g[37], 	p[37], 	x[37]) ;
    _gpx _gpx_38	(a[38],	b[38],	g[38], 	p[38], 	x[38]) ;
    _gpx _gpx_39	(a[39],	b[39],	g[39], 	p[39], 	x[39]) ;
    _gpx _gpx_40	(a[40],	b[40],	g[40], 	p[40], 	x[40]) ;
    _gpx _gpx_41	(a[41],	b[41],	g[41], 	p[41], 	x[41]) ;
    _gpx _gpx_42	(a[42],	b[42],	g[42], 	p[42], 	x[42]) ;
    _gpx _gpx_43	(a[43],	b[43],	g[43], 	p[43], 	x[43]) ;
    _gpx _gpx_44	(a[44],	b[44],	g[44], 	p[44], 	x[44]) ;
    _gpx _gpx_45	(a[45],	b[45],	g[45], 	p[45], 	x[45]) ;
    _gpx _gpx_46	(a[46],	b[46],	g[46], 	p[46], 	x[46]) ;
    _gpx _gpx_47	(a[47],	b[47],	g[47], 	p[47], 	x[47]) ;
    _gpx _gpx_48	(a[48],	b[48],	g[48], 	p[48], 	x[48]) ;
    _gpx _gpx_49	(a[49],	b[49],	g[49], 	p[49], 	x[49]) ;
    _gpx _gpx_50	(a[50],	b[50],	g[50], 	p[50], 	x[50]) ;
    _gpx _gpx_51	(a[51],	b[51],	g[51], 	p[51], 	x[51]) ;
    _gpx _gpx_52	(a[52],	b[52],	g[52], 	p[52], 	x[52]) ;
    _gpx _gpx_53	(a[53],	b[53],	g[53], 	p[53], 	x[53]) ;
    _gpx _gpx_54	(a[54],	b[54],	g[54], 	p[54], 	x[54]) ;
    _gpx _gpx_55	(a[55],	b[55],	g[55], 	p[55], 	x[55]) ;
    _gpx _gpx_56	(a[56],	b[56],	g[56], 	p[56], 	x[56]) ;
    _gpx _gpx_57	(a[57],	b[57],	g[57], 	p[57], 	x[57]) ;
    _gpx _gpx_58	(a[58],	b[58],	g[58], 	p[58], 	x[58]) ;
    _gpx _gpx_59	(a[59],	b[59],	g[59], 	p[59], 	x[59]) ;
    _gpx _gpx_60	(a[60],	b[60],	g[60], 	p[60], 	x[60]) ;
    _gpx _gpx_61	(a[61],	b[61],	g[61], 	p[61], 	x[61]) ;
    _gpx _gpx_62	(a[62],	b[62],	g[62], 	p[62], 	x[62]) ;
    _gpx _gpx_63	(a[63],	b[63],	g[63], 	p[63], 	x[63]) ;

    _4g2p_H4 _4g2p_H4_0( {g[0],g[63],g[62],g[61]} ,{p[63],p[62]} , H1[0] ) ;
    _4g2p_H4 _4g2p_H4_1( {g[1],g[0],g[63],g[62]} ,{p[0],p[63]} , H1[1] ) ;
    _4g2p_H4 _4g2p_H4_2( {g[2],g[1],g[0],g[63]} ,{p[1],p[0]} , H1[2] ) ;
    _4g2p_H4 _4g2p_H4_3( {g[3],g[2],g[1],g[0]} ,{p[2],p[1]} , H1[3] ) ;
    _4g2p_H4 _4g2p_H4_4( {g[4],g[3],g[2],g[1]} ,{p[3],p[2]} , H1[4] ) ;
    _4g2p_H4 _4g2p_H4_5( {g[5],g[4],g[3],g[2]} ,{p[4],p[3]} , H1[5] ) ;
    _4g2p_H4 _4g2p_H4_6( {g[6],g[5],g[4],g[3]} ,{p[5],p[4]} , H1[6] ) ;
    _4g2p_H4 _4g2p_H4_7( {g[7],g[6],g[5],g[4]} ,{p[6],p[5]} , H1[7] ) ;
    _4g2p_H4 _4g2p_H4_8( {g[8],g[7],g[6],g[5]} ,{p[7],p[6]} , H1[8] ) ;
    _4g2p_H4 _4g2p_H4_9( {g[9],g[8],g[7],g[6]} ,{p[8],p[7]} , H1[9] ) ;
    _4g2p_H4 _4g2p_H4_10( {g[10],g[9],g[8],g[7]} ,{p[9],p[8]} , H1[10] ) ;
    _4g2p_H4 _4g2p_H4_11( {g[11],g[10],g[9],g[8]} ,{p[10],p[9]} , H1[11] ) ;
    _4g2p_H4 _4g2p_H4_12( {g[12],g[11],g[10],g[9]} ,{p[11],p[10]} , H1[12] ) ;
    _4g2p_H4 _4g2p_H4_13( {g[13],g[12],g[11],g[10]} ,{p[12],p[11]} , H1[13] ) ;
    _4g2p_H4 _4g2p_H4_14( {g[14],g[13],g[12],g[11]} ,{p[13],p[12]} , H1[14] ) ;
    _4g2p_H4 _4g2p_H4_15( {g[15],g[14],g[13],g[12]} ,{p[14],p[13]} , H1[15] ) ;
    _4g2p_H4 _4g2p_H4_16( {g[16],g[15],g[14],g[13]} ,{p[15],p[14]} , H1[16] ) ;
    _4g2p_H4 _4g2p_H4_17( {g[17],g[16],g[15],g[14]} ,{p[16],p[15]} , H1[17] ) ;
    _4g2p_H4 _4g2p_H4_18( {g[18],g[17],g[16],g[15]} ,{p[17],p[16]} , H1[18] ) ;
    _4g2p_H4 _4g2p_H4_19( {g[19],g[18],g[17],g[16]} ,{p[18],p[17]} , H1[19] ) ;
    _4g2p_H4 _4g2p_H4_20( {g[20],g[19],g[18],g[17]} ,{p[19],p[18]} , H1[20] ) ;
    _4g2p_H4 _4g2p_H4_21( {g[21],g[20],g[19],g[18]} ,{p[20],p[19]} , H1[21] ) ;
    _4g2p_H4 _4g2p_H4_22( {g[22],g[21],g[20],g[19]} ,{p[21],p[20]} , H1[22] ) ;
    _4g2p_H4 _4g2p_H4_23( {g[23],g[22],g[21],g[20]} ,{p[22],p[21]} , H1[23] ) ;
    _4g2p_H4 _4g2p_H4_24( {g[24],g[23],g[22],g[21]} ,{p[23],p[22]} , H1[24] ) ;
    _4g2p_H4 _4g2p_H4_25( {g[25],g[24],g[23],g[22]} ,{p[24],p[23]} , H1[25] ) ;
    _4g2p_H4 _4g2p_H4_26( {g[26],g[25],g[24],g[23]} ,{p[25],p[24]} , H1[26] ) ;
    _4g2p_H4 _4g2p_H4_27( {g[27],g[26],g[25],g[24]} ,{p[26],p[25]} , H1[27] ) ;
    _4g2p_H4 _4g2p_H4_28( {g[28],g[27],g[26],g[25]} ,{p[27],p[26]} , H1[28] ) ;
    _4g2p_H4 _4g2p_H4_29( {g[29],g[28],g[27],g[26]} ,{p[28],p[27]} , H1[29] ) ;
    _4g2p_H4 _4g2p_H4_30( {g[30],g[29],g[28],g[27]} ,{p[29],p[28]} , H1[30] ) ;
    _4g2p_H4 _4g2p_H4_31( {g[31],g[30],g[29],g[28]} ,{p[30],p[29]} , H1[31] ) ;
    _4g2p_H4 _4g2p_H4_32( {g[32],g[31],g[30],g[29]} ,{p[31],p[30]} , H1[32] ) ;
    _4g2p_H4 _4g2p_H4_33( {g[33],g[32],g[31],g[30]} ,{p[32],p[31]} , H1[33] ) ;
    _4g2p_H4 _4g2p_H4_34( {g[34],g[33],g[32],g[31]} ,{p[33],p[32]} , H1[34] ) ;
    _4g2p_H4 _4g2p_H4_35( {g[35],g[34],g[33],g[32]} ,{p[34],p[33]} , H1[35] ) ;
    _4g2p_H4 _4g2p_H4_36( {g[36],g[35],g[34],g[33]} ,{p[35],p[34]} , H1[36] ) ;
    _4g2p_H4 _4g2p_H4_37( {g[37],g[36],g[35],g[34]} ,{p[36],p[35]} , H1[37] ) ;
    _4g2p_H4 _4g2p_H4_38( {g[38],g[37],g[36],g[35]} ,{p[37],p[36]} , H1[38] ) ;
    _4g2p_H4 _4g2p_H4_39( {g[39],g[38],g[37],g[36]} ,{p[38],p[37]} , H1[39] ) ;
    _4g2p_H4 _4g2p_H4_40( {g[40],g[39],g[38],g[37]} ,{p[39],p[38]} , H1[40] ) ;
    _4g2p_H4 _4g2p_H4_41( {g[41],g[40],g[39],g[38]} ,{p[40],p[39]} , H1[41] ) ;
    _4g2p_H4 _4g2p_H4_42( {g[42],g[41],g[40],g[39]} ,{p[41],p[40]} , H1[42] ) ;
    _4g2p_H4 _4g2p_H4_43( {g[43],g[42],g[41],g[40]} ,{p[42],p[41]} , H1[43] ) ;
    _4g2p_H4 _4g2p_H4_44( {g[44],g[43],g[42],g[41]} ,{p[43],p[42]} , H1[44] ) ;
    _4g2p_H4 _4g2p_H4_45( {g[45],g[44],g[43],g[42]} ,{p[44],p[43]} , H1[45] ) ;
    _4g2p_H4 _4g2p_H4_46( {g[46],g[45],g[44],g[43]} ,{p[45],p[44]} , H1[46] ) ;
    _4g2p_H4 _4g2p_H4_47( {g[47],g[46],g[45],g[44]} ,{p[46],p[45]} , H1[47] ) ;
    _4g2p_H4 _4g2p_H4_48( {g[48],g[47],g[46],g[45]} ,{p[47],p[46]} , H1[48] ) ;
    _4g2p_H4 _4g2p_H4_49( {g[49],g[48],g[47],g[46]} ,{p[48],p[47]} , H1[49] ) ;
    _4g2p_H4 _4g2p_H4_50( {g[50],g[49],g[48],g[47]} ,{p[49],p[48]} , H1[50] ) ;
    _4g2p_H4 _4g2p_H4_51( {g[51],g[50],g[49],g[48]} ,{p[50],p[49]} , H1[51] ) ;
    _4g2p_H4 _4g2p_H4_52( {g[52],g[51],g[50],g[49]} ,{p[51],p[50]} , H1[52] ) ;
    _4g2p_H4 _4g2p_H4_53( {g[53],g[52],g[51],g[50]} ,{p[52],p[51]} , H1[53] ) ;
    _4g2p_H4 _4g2p_H4_54( {g[54],g[53],g[52],g[51]} ,{p[53],p[52]} , H1[54] ) ;
    _4g2p_H4 _4g2p_H4_55( {g[55],g[54],g[53],g[52]} ,{p[54],p[53]} , H1[55] ) ;
    _4g2p_H4 _4g2p_H4_56( {g[56],g[55],g[54],g[53]} ,{p[55],p[54]} , H1[56] ) ;
    _4g2p_H4 _4g2p_H4_57( {g[57],g[56],g[55],g[54]} ,{p[56],p[55]} , H1[57] ) ;
    _4g2p_H4 _4g2p_H4_58( {g[58],g[57],g[56],g[55]} ,{p[57],p[56]} , H1[58] ) ;
    _4g2p_H4 _4g2p_H4_59( {g[59],g[58],g[57],g[56]} ,{p[58],p[57]} , H1[59] ) ;
    _4g2p_H4 _4g2p_H4_60( {g[60],g[59],g[58],g[57]} ,{p[59],p[58]} , H1[60] ) ;
    _4g2p_H4 _4g2p_H4_61( {g[61],g[60],g[59],g[58]} ,{p[60],p[59]} , H1[61] ) ;
    _4g2p_H4 _4g2p_H4_62( {g[62],g[61],g[60],g[59]} ,{p[61],p[60]} , H1[62] ) ;
    _4g2p_H4 _4g2p_H4_63( {g[63],g[62],g[61],g[60]} ,{p[62],p[61]} , H1[63] ) ;

    _P4 _P4_0( {p[0],p[63],p[62],p[61]} ,Pr1[0] ) ;
    _P4 _P4_1( {p[1],p[0],p[63],p[62]} ,Pr1[1] ) ;
    _P4 _P4_2( {p[2],p[1],p[0],p[63]} ,Pr1[2] ) ;
    _P4 _P4_3( {p[3],p[2],p[1],p[0]} ,Pr1[3] ) ;
    _P4 _P4_4( {p[4],p[3],p[2],p[1]} ,Pr1[4] ) ;
    _P4 _P4_5( {p[5],p[4],p[3],p[2]} ,Pr1[5] ) ;
    _P4 _P4_6( {p[6],p[5],p[4],p[3]} ,Pr1[6] ) ;
    _P4 _P4_7( {p[7],p[6],p[5],p[4]} ,Pr1[7] ) ;
    _P4 _P4_8( {p[8],p[7],p[6],p[5]} ,Pr1[8] ) ;
    _P4 _P4_9( {p[9],p[8],p[7],p[6]} ,Pr1[9] ) ;
    _P4 _P4_10( {p[10],p[9],p[8],p[7]} ,Pr1[10] ) ;
    _P4 _P4_11( {p[11],p[10],p[9],p[8]} ,Pr1[11] ) ;
    _P4 _P4_12( {p[12],p[11],p[10],p[9]} ,Pr1[12] ) ;
    _P4 _P4_13( {p[13],p[12],p[11],p[10]} ,Pr1[13] ) ;
    _P4 _P4_14( {p[14],p[13],p[12],p[11]} ,Pr1[14] ) ;
    _P4 _P4_15( {p[15],p[14],p[13],p[12]} ,Pr1[15] ) ;
    _P4 _P4_16( {p[16],p[15],p[14],p[13]} ,Pr1[16] ) ;
    _P4 _P4_17( {p[17],p[16],p[15],p[14]} ,Pr1[17] ) ;
    _P4 _P4_18( {p[18],p[17],p[16],p[15]} ,Pr1[18] ) ;
    _P4 _P4_19( {p[19],p[18],p[17],p[16]} ,Pr1[19] ) ;
    _P4 _P4_20( {p[20],p[19],p[18],p[17]} ,Pr1[20] ) ;
    _P4 _P4_21( {p[21],p[20],p[19],p[18]} ,Pr1[21] ) ;
    _P4 _P4_22( {p[22],p[21],p[20],p[19]} ,Pr1[22] ) ;
    _P4 _P4_23( {p[23],p[22],p[21],p[20]} ,Pr1[23] ) ;
    _P4 _P4_24( {p[24],p[23],p[22],p[21]} ,Pr1[24] ) ;
    _P4 _P4_25( {p[25],p[24],p[23],p[22]} ,Pr1[25] ) ;
    _P4 _P4_26( {p[26],p[25],p[24],p[23]} ,Pr1[26] ) ;
    _P4 _P4_27( {p[27],p[26],p[25],p[24]} ,Pr1[27] ) ;
    _P4 _P4_28( {p[28],p[27],p[26],p[25]} ,Pr1[28] ) ;
    _P4 _P4_29( {p[29],p[28],p[27],p[26]} ,Pr1[29] ) ;
    _P4 _P4_30( {p[30],p[29],p[28],p[27]} ,Pr1[30] ) ;
    _P4 _P4_31( {p[31],p[30],p[29],p[28]} ,Pr1[31] ) ;
    _P4 _P4_32( {p[32],p[31],p[30],p[29]} ,Pr1[32] ) ;
    _P4 _P4_33( {p[33],p[32],p[31],p[30]} ,Pr1[33] ) ;
    _P4 _P4_34( {p[34],p[33],p[32],p[31]} ,Pr1[34] ) ;
    _P4 _P4_35( {p[35],p[34],p[33],p[32]} ,Pr1[35] ) ;
    _P4 _P4_36( {p[36],p[35],p[34],p[33]} ,Pr1[36] ) ;
    _P4 _P4_37( {p[37],p[36],p[35],p[34]} ,Pr1[37] ) ;
    _P4 _P4_38( {p[38],p[37],p[36],p[35]} ,Pr1[38] ) ;
    _P4 _P4_39( {p[39],p[38],p[37],p[36]} ,Pr1[39] ) ;
    _P4 _P4_40( {p[40],p[39],p[38],p[37]} ,Pr1[40] ) ;
    _P4 _P4_41( {p[41],p[40],p[39],p[38]} ,Pr1[41] ) ;
    _P4 _P4_42( {p[42],p[41],p[40],p[39]} ,Pr1[42] ) ;
    _P4 _P4_43( {p[43],p[42],p[41],p[40]} ,Pr1[43] ) ;
    _P4 _P4_44( {p[44],p[43],p[42],p[41]} ,Pr1[44] ) ;
    _P4 _P4_45( {p[45],p[44],p[43],p[42]} ,Pr1[45] ) ;
    _P4 _P4_46( {p[46],p[45],p[44],p[43]} ,Pr1[46] ) ;
    _P4 _P4_47( {p[47],p[46],p[45],p[44]} ,Pr1[47] ) ;
    _P4 _P4_48( {p[48],p[47],p[46],p[45]} ,Pr1[48] ) ;
    _P4 _P4_49( {p[49],p[48],p[47],p[46]} ,Pr1[49] ) ;
    _P4 _P4_50( {p[50],p[49],p[48],p[47]} ,Pr1[50] ) ;
    _P4 _P4_51( {p[51],p[50],p[49],p[48]} ,Pr1[51] ) ;
    _P4 _P4_52( {p[52],p[51],p[50],p[49]} ,Pr1[52] ) ;
    _P4 _P4_53( {p[53],p[52],p[51],p[50]} ,Pr1[53] ) ;
    _P4 _P4_54( {p[54],p[53],p[52],p[51]} ,Pr1[54] ) ;
    _P4 _P4_55( {p[55],p[54],p[53],p[52]} ,Pr1[55] ) ;
    _P4 _P4_56( {p[56],p[55],p[54],p[53]} ,Pr1[56] ) ;
    _P4 _P4_57( {p[57],p[56],p[55],p[54]} ,Pr1[57] ) ;
    _P4 _P4_58( {p[58],p[57],p[56],p[55]} ,Pr1[58] ) ;
    _P4 _P4_59( {p[59],p[58],p[57],p[56]} ,Pr1[59] ) ;
    _P4 _P4_60( {p[60],p[59],p[58],p[57]} ,Pr1[60] ) ;
    _P4 _P4_61( {p[61],p[60],p[59],p[58]} ,Pr1[61] ) ;
    _P4 _P4_62( {p[62],p[61],p[60],p[59]} ,Pr1[62] ) ;
    _P4 _P4_63( {p[63],p[62],p[61],p[60]} ,Pr1[63] ) ;

    _4G3P_G4 _4G3P_G4_0( {H1[0],H1[60],H1[56],H1[52]} , {Pr1[63],Pr1[59],Pr1[55]} ,H2[0] ) ;
    _4G3P_G4 _4G3P_G4_1( {H1[1],H1[61],H1[57],H1[53]} , {Pr1[0],Pr1[60],Pr1[56]} ,H2[1] ) ;
    _4G3P_G4 _4G3P_G4_2( {H1[2],H1[62],H1[58],H1[54]} , {Pr1[1],Pr1[61],Pr1[57]} ,H2[2] ) ;
    _4G3P_G4 _4G3P_G4_3( {H1[3],H1[63],H1[59],H1[55]} , {Pr1[2],Pr1[62],Pr1[58]} ,H2[3] ) ;
    _4G3P_G4 _4G3P_G4_4( {H1[4],H1[0],H1[60],H1[56]} , {Pr1[3],Pr1[63],Pr1[59]} ,H2[4] ) ;
    _4G3P_G4 _4G3P_G4_5( {H1[5],H1[1],H1[61],H1[57]} , {Pr1[4],Pr1[0],Pr1[60]} ,H2[5] ) ;
    _4G3P_G4 _4G3P_G4_6( {H1[6],H1[2],H1[62],H1[58]} , {Pr1[5],Pr1[1],Pr1[61]} ,H2[6] ) ;
    _4G3P_G4 _4G3P_G4_7( {H1[7],H1[3],H1[63],H1[59]} , {Pr1[6],Pr1[2],Pr1[62]} ,H2[7] ) ;
    _4G3P_G4 _4G3P_G4_8( {H1[8],H1[4],H1[0],H1[60]} , {Pr1[7],Pr1[3],Pr1[63]} ,H2[8] ) ;
    _4G3P_G4 _4G3P_G4_9( {H1[9],H1[5],H1[1],H1[61]} , {Pr1[8],Pr1[4],Pr1[0]} ,H2[9] ) ;
    _4G3P_G4 _4G3P_G4_10( {H1[10],H1[6],H1[2],H1[62]} , {Pr1[9],Pr1[5],Pr1[1]} ,H2[10] ) ;
    _4G3P_G4 _4G3P_G4_11( {H1[11],H1[7],H1[3],H1[63]} , {Pr1[10],Pr1[6],Pr1[2]} ,H2[11] ) ;
    _4G3P_G4 _4G3P_G4_12( {H1[12],H1[8],H1[4],H1[0]} , {Pr1[11],Pr1[7],Pr1[3]} ,H2[12] ) ;
    _4G3P_G4 _4G3P_G4_13( {H1[13],H1[9],H1[5],H1[1]} , {Pr1[12],Pr1[8],Pr1[4]} ,H2[13] ) ;
    _4G3P_G4 _4G3P_G4_14( {H1[14],H1[10],H1[6],H1[2]} , {Pr1[13],Pr1[9],Pr1[5]} ,H2[14] ) ;
    _4G3P_G4 _4G3P_G4_15( {H1[15],H1[11],H1[7],H1[3]} , {Pr1[14],Pr1[10],Pr1[6]} ,H2[15] ) ;
    _4G3P_G4 _4G3P_G4_16( {H1[16],H1[12],H1[8],H1[4]} , {Pr1[15],Pr1[11],Pr1[7]} ,H2[16] ) ;
    _4G3P_G4 _4G3P_G4_17( {H1[17],H1[13],H1[9],H1[5]} , {Pr1[16],Pr1[12],Pr1[8]} ,H2[17] ) ;
    _4G3P_G4 _4G3P_G4_18( {H1[18],H1[14],H1[10],H1[6]} , {Pr1[17],Pr1[13],Pr1[9]} ,H2[18] ) ;
    _4G3P_G4 _4G3P_G4_19( {H1[19],H1[15],H1[11],H1[7]} , {Pr1[18],Pr1[14],Pr1[10]} ,H2[19] ) ;
    _4G3P_G4 _4G3P_G4_20( {H1[20],H1[16],H1[12],H1[8]} , {Pr1[19],Pr1[15],Pr1[11]} ,H2[20] ) ;
    _4G3P_G4 _4G3P_G4_21( {H1[21],H1[17],H1[13],H1[9]} , {Pr1[20],Pr1[16],Pr1[12]} ,H2[21] ) ;
    _4G3P_G4 _4G3P_G4_22( {H1[22],H1[18],H1[14],H1[10]} , {Pr1[21],Pr1[17],Pr1[13]} ,H2[22] ) ;
    _4G3P_G4 _4G3P_G4_23( {H1[23],H1[19],H1[15],H1[11]} , {Pr1[22],Pr1[18],Pr1[14]} ,H2[23] ) ;
    _4G3P_G4 _4G3P_G4_24( {H1[24],H1[20],H1[16],H1[12]} , {Pr1[23],Pr1[19],Pr1[15]} ,H2[24] ) ;
    _4G3P_G4 _4G3P_G4_25( {H1[25],H1[21],H1[17],H1[13]} , {Pr1[24],Pr1[20],Pr1[16]} ,H2[25] ) ;
    _4G3P_G4 _4G3P_G4_26( {H1[26],H1[22],H1[18],H1[14]} , {Pr1[25],Pr1[21],Pr1[17]} ,H2[26] ) ;
    _4G3P_G4 _4G3P_G4_27( {H1[27],H1[23],H1[19],H1[15]} , {Pr1[26],Pr1[22],Pr1[18]} ,H2[27] ) ;
    _4G3P_G4 _4G3P_G4_28( {H1[28],H1[24],H1[20],H1[16]} , {Pr1[27],Pr1[23],Pr1[19]} ,H2[28] ) ;
    _4G3P_G4 _4G3P_G4_29( {H1[29],H1[25],H1[21],H1[17]} , {Pr1[28],Pr1[24],Pr1[20]} ,H2[29] ) ;
    _4G3P_G4 _4G3P_G4_30( {H1[30],H1[26],H1[22],H1[18]} , {Pr1[29],Pr1[25],Pr1[21]} ,H2[30] ) ;
    _4G3P_G4 _4G3P_G4_31( {H1[31],H1[27],H1[23],H1[19]} , {Pr1[30],Pr1[26],Pr1[22]} ,H2[31] ) ;
    _4G3P_G4 _4G3P_G4_32( {H1[32],H1[28],H1[24],H1[20]} , {Pr1[31],Pr1[27],Pr1[23]} ,H2[32] ) ;
    _4G3P_G4 _4G3P_G4_33( {H1[33],H1[29],H1[25],H1[21]} , {Pr1[32],Pr1[28],Pr1[24]} ,H2[33] ) ;
    _4G3P_G4 _4G3P_G4_34( {H1[34],H1[30],H1[26],H1[22]} , {Pr1[33],Pr1[29],Pr1[25]} ,H2[34] ) ;
    _4G3P_G4 _4G3P_G4_35( {H1[35],H1[31],H1[27],H1[23]} , {Pr1[34],Pr1[30],Pr1[26]} ,H2[35] ) ;
    _4G3P_G4 _4G3P_G4_36( {H1[36],H1[32],H1[28],H1[24]} , {Pr1[35],Pr1[31],Pr1[27]} ,H2[36] ) ;
    _4G3P_G4 _4G3P_G4_37( {H1[37],H1[33],H1[29],H1[25]} , {Pr1[36],Pr1[32],Pr1[28]} ,H2[37] ) ;
    _4G3P_G4 _4G3P_G4_38( {H1[38],H1[34],H1[30],H1[26]} , {Pr1[37],Pr1[33],Pr1[29]} ,H2[38] ) ;
    _4G3P_G4 _4G3P_G4_39( {H1[39],H1[35],H1[31],H1[27]} , {Pr1[38],Pr1[34],Pr1[30]} ,H2[39] ) ;
    _4G3P_G4 _4G3P_G4_40( {H1[40],H1[36],H1[32],H1[28]} , {Pr1[39],Pr1[35],Pr1[31]} ,H2[40] ) ;
    _4G3P_G4 _4G3P_G4_41( {H1[41],H1[37],H1[33],H1[29]} , {Pr1[40],Pr1[36],Pr1[32]} ,H2[41] ) ;
    _4G3P_G4 _4G3P_G4_42( {H1[42],H1[38],H1[34],H1[30]} , {Pr1[41],Pr1[37],Pr1[33]} ,H2[42] ) ;
    _4G3P_G4 _4G3P_G4_43( {H1[43],H1[39],H1[35],H1[31]} , {Pr1[42],Pr1[38],Pr1[34]} ,H2[43] ) ;
    _4G3P_G4 _4G3P_G4_44( {H1[44],H1[40],H1[36],H1[32]} , {Pr1[43],Pr1[39],Pr1[35]} ,H2[44] ) ;
    _4G3P_G4 _4G3P_G4_45( {H1[45],H1[41],H1[37],H1[33]} , {Pr1[44],Pr1[40],Pr1[36]} ,H2[45] ) ;
    _4G3P_G4 _4G3P_G4_46( {H1[46],H1[42],H1[38],H1[34]} , {Pr1[45],Pr1[41],Pr1[37]} ,H2[46] ) ;
    _4G3P_G4 _4G3P_G4_47( {H1[47],H1[43],H1[39],H1[35]} , {Pr1[46],Pr1[42],Pr1[38]} ,H2[47] ) ;
    _4G3P_G4 _4G3P_G4_48( {H1[48],H1[44],H1[40],H1[36]} , {Pr1[47],Pr1[43],Pr1[39]} ,H2[48] ) ;
    _4G3P_G4 _4G3P_G4_49( {H1[49],H1[45],H1[41],H1[37]} , {Pr1[48],Pr1[44],Pr1[40]} ,H2[49] ) ;
    _4G3P_G4 _4G3P_G4_50( {H1[50],H1[46],H1[42],H1[38]} , {Pr1[49],Pr1[45],Pr1[41]} ,H2[50] ) ;
    _4G3P_G4 _4G3P_G4_51( {H1[51],H1[47],H1[43],H1[39]} , {Pr1[50],Pr1[46],Pr1[42]} ,H2[51] ) ;
    _4G3P_G4 _4G3P_G4_52( {H1[52],H1[48],H1[44],H1[40]} , {Pr1[51],Pr1[47],Pr1[43]} ,H2[52] ) ;
    _4G3P_G4 _4G3P_G4_53( {H1[53],H1[49],H1[45],H1[41]} , {Pr1[52],Pr1[48],Pr1[44]} ,H2[53] ) ;
    _4G3P_G4 _4G3P_G4_54( {H1[54],H1[50],H1[46],H1[42]} , {Pr1[53],Pr1[49],Pr1[45]} ,H2[54] ) ;
    _4G3P_G4 _4G3P_G4_55( {H1[55],H1[51],H1[47],H1[43]} , {Pr1[54],Pr1[50],Pr1[46]} ,H2[55] ) ;
    _4G3P_G4 _4G3P_G4_56( {H1[56],H1[52],H1[48],H1[44]} , {Pr1[55],Pr1[51],Pr1[47]} ,H2[56] ) ;
    _4G3P_G4 _4G3P_G4_57( {H1[57],H1[53],H1[49],H1[45]} , {Pr1[56],Pr1[52],Pr1[48]} ,H2[57] ) ;
    _4G3P_G4 _4G3P_G4_58( {H1[58],H1[54],H1[50],H1[46]} , {Pr1[57],Pr1[53],Pr1[49]} ,H2[58] ) ;
    _4G3P_G4 _4G3P_G4_59( {H1[59],H1[55],H1[51],H1[47]} , {Pr1[58],Pr1[54],Pr1[50]} ,H2[59] ) ;
    _4G3P_G4 _4G3P_G4_60( {H1[60],H1[56],H1[52],H1[48]} , {Pr1[59],Pr1[55],Pr1[51]} ,H2[60] ) ;
    _4G3P_G4 _4G3P_G4_61( {H1[61],H1[57],H1[53],H1[49]} , {Pr1[60],Pr1[56],Pr1[52]} ,H2[61] ) ;
    _4G3P_G4 _4G3P_G4_62( {H1[62],H1[58],H1[54],H1[50]} , {Pr1[61],Pr1[57],Pr1[53]} ,H2[62] ) ;
    _4G3P_G4 _4G3P_G4_63( {H1[63],H1[59],H1[55],H1[51]} , {Pr1[62],Pr1[58],Pr1[54]} ,H2[63] ) ;

    _P4 _P4_64( {Pr1[0],Pr1[60],Pr1[56],Pr1[52]} ,Pr2[0] ) ;
    _P4 _P4_65( {Pr1[1],Pr1[61],Pr1[57],Pr1[53]} ,Pr2[1] ) ;
    _P4 _P4_66( {Pr1[2],Pr1[62],Pr1[58],Pr1[54]} ,Pr2[2] ) ;
    _P4 _P4_67( {Pr1[3],Pr1[63],Pr1[59],Pr1[55]} ,Pr2[3] ) ;
    _P4 _P4_68( {Pr1[4],Pr1[0],Pr1[60],Pr1[56]} ,Pr2[4] ) ;
    _P4 _P4_69( {Pr1[5],Pr1[1],Pr1[61],Pr1[57]} ,Pr2[5] ) ;
    _P4 _P4_70( {Pr1[6],Pr1[2],Pr1[62],Pr1[58]} ,Pr2[6] ) ;
    _P4 _P4_71( {Pr1[7],Pr1[3],Pr1[63],Pr1[59]} ,Pr2[7] ) ;
    _P4 _P4_72( {Pr1[8],Pr1[4],Pr1[0],Pr1[60]} ,Pr2[8] ) ;
    _P4 _P4_73( {Pr1[9],Pr1[5],Pr1[1],Pr1[61]} ,Pr2[9] ) ;
    _P4 _P4_74( {Pr1[10],Pr1[6],Pr1[2],Pr1[62]} ,Pr2[10] ) ;
    _P4 _P4_75( {Pr1[11],Pr1[7],Pr1[3],Pr1[63]} ,Pr2[11] ) ;
    _P4 _P4_76( {Pr1[12],Pr1[8],Pr1[4],Pr1[0]} ,Pr2[12] ) ;
    _P4 _P4_77( {Pr1[13],Pr1[9],Pr1[5],Pr1[1]} ,Pr2[13] ) ;
    _P4 _P4_78( {Pr1[14],Pr1[10],Pr1[6],Pr1[2]} ,Pr2[14] ) ;
    _P4 _P4_79( {Pr1[15],Pr1[11],Pr1[7],Pr1[3]} ,Pr2[15] ) ;
    _P4 _P4_80( {Pr1[16],Pr1[12],Pr1[8],Pr1[4]} ,Pr2[16] ) ;
    _P4 _P4_81( {Pr1[17],Pr1[13],Pr1[9],Pr1[5]} ,Pr2[17] ) ;
    _P4 _P4_82( {Pr1[18],Pr1[14],Pr1[10],Pr1[6]} ,Pr2[18] ) ;
    _P4 _P4_83( {Pr1[19],Pr1[15],Pr1[11],Pr1[7]} ,Pr2[19] ) ;
    _P4 _P4_84( {Pr1[20],Pr1[16],Pr1[12],Pr1[8]} ,Pr2[20] ) ;
    _P4 _P4_85( {Pr1[21],Pr1[17],Pr1[13],Pr1[9]} ,Pr2[21] ) ;
    _P4 _P4_86( {Pr1[22],Pr1[18],Pr1[14],Pr1[10]} ,Pr2[22] ) ;
    _P4 _P4_87( {Pr1[23],Pr1[19],Pr1[15],Pr1[11]} ,Pr2[23] ) ;
    _P4 _P4_88( {Pr1[24],Pr1[20],Pr1[16],Pr1[12]} ,Pr2[24] ) ;
    _P4 _P4_89( {Pr1[25],Pr1[21],Pr1[17],Pr1[13]} ,Pr2[25] ) ;
    _P4 _P4_90( {Pr1[26],Pr1[22],Pr1[18],Pr1[14]} ,Pr2[26] ) ;
    _P4 _P4_91( {Pr1[27],Pr1[23],Pr1[19],Pr1[15]} ,Pr2[27] ) ;
    _P4 _P4_92( {Pr1[28],Pr1[24],Pr1[20],Pr1[16]} ,Pr2[28] ) ;
    _P4 _P4_93( {Pr1[29],Pr1[25],Pr1[21],Pr1[17]} ,Pr2[29] ) ;
    _P4 _P4_94( {Pr1[30],Pr1[26],Pr1[22],Pr1[18]} ,Pr2[30] ) ;
    _P4 _P4_95( {Pr1[31],Pr1[27],Pr1[23],Pr1[19]} ,Pr2[31] ) ;
    _P4 _P4_96( {Pr1[32],Pr1[28],Pr1[24],Pr1[20]} ,Pr2[32] ) ;
    _P4 _P4_97( {Pr1[33],Pr1[29],Pr1[25],Pr1[21]} ,Pr2[33] ) ;
    _P4 _P4_98( {Pr1[34],Pr1[30],Pr1[26],Pr1[22]} ,Pr2[34] ) ;
    _P4 _P4_99( {Pr1[35],Pr1[31],Pr1[27],Pr1[23]} ,Pr2[35] ) ;
    _P4 _P4_100( {Pr1[36],Pr1[32],Pr1[28],Pr1[24]} ,Pr2[36] ) ;
    _P4 _P4_101( {Pr1[37],Pr1[33],Pr1[29],Pr1[25]} ,Pr2[37] ) ;
    _P4 _P4_102( {Pr1[38],Pr1[34],Pr1[30],Pr1[26]} ,Pr2[38] ) ;
    _P4 _P4_103( {Pr1[39],Pr1[35],Pr1[31],Pr1[27]} ,Pr2[39] ) ;
    _P4 _P4_104( {Pr1[40],Pr1[36],Pr1[32],Pr1[28]} ,Pr2[40] ) ;
    _P4 _P4_105( {Pr1[41],Pr1[37],Pr1[33],Pr1[29]} ,Pr2[41] ) ;
    _P4 _P4_106( {Pr1[42],Pr1[38],Pr1[34],Pr1[30]} ,Pr2[42] ) ;
    _P4 _P4_107( {Pr1[43],Pr1[39],Pr1[35],Pr1[31]} ,Pr2[43] ) ;
    _P4 _P4_108( {Pr1[44],Pr1[40],Pr1[36],Pr1[32]} ,Pr2[44] ) ;
    _P4 _P4_109( {Pr1[45],Pr1[41],Pr1[37],Pr1[33]} ,Pr2[45] ) ;
    _P4 _P4_110( {Pr1[46],Pr1[42],Pr1[38],Pr1[34]} ,Pr2[46] ) ;
    _P4 _P4_111( {Pr1[47],Pr1[43],Pr1[39],Pr1[35]} ,Pr2[47] ) ;
    _P4 _P4_112( {Pr1[48],Pr1[44],Pr1[40],Pr1[36]} ,Pr2[48] ) ;
    _P4 _P4_113( {Pr1[49],Pr1[45],Pr1[41],Pr1[37]} ,Pr2[49] ) ;
    _P4 _P4_114( {Pr1[50],Pr1[46],Pr1[42],Pr1[38]} ,Pr2[50] ) ;
    _P4 _P4_115( {Pr1[51],Pr1[47],Pr1[43],Pr1[39]} ,Pr2[51] ) ;
    _P4 _P4_116( {Pr1[52],Pr1[48],Pr1[44],Pr1[40]} ,Pr2[52] ) ;
    _P4 _P4_117( {Pr1[53],Pr1[49],Pr1[45],Pr1[41]} ,Pr2[53] ) ;
    _P4 _P4_118( {Pr1[54],Pr1[50],Pr1[46],Pr1[42]} ,Pr2[54] ) ;
    _P4 _P4_119( {Pr1[55],Pr1[51],Pr1[47],Pr1[43]} ,Pr2[55] ) ;
    _P4 _P4_120( {Pr1[56],Pr1[52],Pr1[48],Pr1[44]} ,Pr2[56] ) ;
    _P4 _P4_121( {Pr1[57],Pr1[53],Pr1[49],Pr1[45]} ,Pr2[57] ) ;
    _P4 _P4_122( {Pr1[58],Pr1[54],Pr1[50],Pr1[46]} ,Pr2[58] ) ;
    _P4 _P4_123( {Pr1[59],Pr1[55],Pr1[51],Pr1[47]} ,Pr2[59] ) ;
    _P4 _P4_124( {Pr1[60],Pr1[56],Pr1[52],Pr1[48]} ,Pr2[60] ) ;
    _P4 _P4_125( {Pr1[61],Pr1[57],Pr1[53],Pr1[49]} ,Pr2[61] ) ;
    _P4 _P4_126( {Pr1[62],Pr1[58],Pr1[54],Pr1[50]} ,Pr2[62] ) ;
    _P4 _P4_127( {Pr1[63],Pr1[59],Pr1[55],Pr1[51]} ,Pr2[63] ) ;

    _4G3P_G4 _4G3P_G4_64( {H2[0],H2[48],H2[32],H2[16]} , {Pr2[63],Pr2[47],Pr2[31]} ,H3[0] ) ;
    _4G3P_G4 _4G3P_G4_65( {H2[1],H2[49],H2[33],H2[17]} , {Pr2[0],Pr2[48],Pr2[32]} ,H3[1] ) ;
    _4G3P_G4 _4G3P_G4_66( {H2[2],H2[50],H2[34],H2[18]} , {Pr2[1],Pr2[49],Pr2[33]} ,H3[2] ) ;
    _4G3P_G4 _4G3P_G4_67( {H2[3],H2[51],H2[35],H2[19]} , {Pr2[2],Pr2[50],Pr2[34]} ,H3[3] ) ;
    _4G3P_G4 _4G3P_G4_68( {H2[4],H2[52],H2[36],H2[20]} , {Pr2[3],Pr2[51],Pr2[35]} ,H3[4] ) ;
    _4G3P_G4 _4G3P_G4_69( {H2[5],H2[53],H2[37],H2[21]} , {Pr2[4],Pr2[52],Pr2[36]} ,H3[5] ) ;
    _4G3P_G4 _4G3P_G4_70( {H2[6],H2[54],H2[38],H2[22]} , {Pr2[5],Pr2[53],Pr2[37]} ,H3[6] ) ;
    _4G3P_G4 _4G3P_G4_71( {H2[7],H2[55],H2[39],H2[23]} , {Pr2[6],Pr2[54],Pr2[38]} ,H3[7] ) ;
    _4G3P_G4 _4G3P_G4_72( {H2[8],H2[56],H2[40],H2[24]} , {Pr2[7],Pr2[55],Pr2[39]} ,H3[8] ) ;
    _4G3P_G4 _4G3P_G4_73( {H2[9],H2[57],H2[41],H2[25]} , {Pr2[8],Pr2[56],Pr2[40]} ,H3[9] ) ;
    _4G3P_G4 _4G3P_G4_74( {H2[10],H2[58],H2[42],H2[26]} , {Pr2[9],Pr2[57],Pr2[41]} ,H3[10] ) ;
    _4G3P_G4 _4G3P_G4_75( {H2[11],H2[59],H2[43],H2[27]} , {Pr2[10],Pr2[58],Pr2[42]} ,H3[11] ) ;
    _4G3P_G4 _4G3P_G4_76( {H2[12],H2[60],H2[44],H2[28]} , {Pr2[11],Pr2[59],Pr2[43]} ,H3[12] ) ;
    _4G3P_G4 _4G3P_G4_77( {H2[13],H2[61],H2[45],H2[29]} , {Pr2[12],Pr2[60],Pr2[44]} ,H3[13] ) ;
    _4G3P_G4 _4G3P_G4_78( {H2[14],H2[62],H2[46],H2[30]} , {Pr2[13],Pr2[61],Pr2[45]} ,H3[14] ) ;
    _4G3P_G4 _4G3P_G4_79( {H2[15],H2[63],H2[47],H2[31]} , {Pr2[14],Pr2[62],Pr2[46]} ,H3[15] ) ;
    _4G3P_G4 _4G3P_G4_80( {H2[16],H2[0],H2[48],H2[32]} , {Pr2[15],Pr2[63],Pr2[47]} ,H3[16] ) ;
    _4G3P_G4 _4G3P_G4_81( {H2[17],H2[1],H2[49],H2[33]} , {Pr2[16],Pr2[0],Pr2[48]} ,H3[17] ) ;
    _4G3P_G4 _4G3P_G4_82( {H2[18],H2[2],H2[50],H2[34]} , {Pr2[17],Pr2[1],Pr2[49]} ,H3[18] ) ;
    _4G3P_G4 _4G3P_G4_83( {H2[19],H2[3],H2[51],H2[35]} , {Pr2[18],Pr2[2],Pr2[50]} ,H3[19] ) ;
    _4G3P_G4 _4G3P_G4_84( {H2[20],H2[4],H2[52],H2[36]} , {Pr2[19],Pr2[3],Pr2[51]} ,H3[20] ) ;
    _4G3P_G4 _4G3P_G4_85( {H2[21],H2[5],H2[53],H2[37]} , {Pr2[20],Pr2[4],Pr2[52]} ,H3[21] ) ;
    _4G3P_G4 _4G3P_G4_86( {H2[22],H2[6],H2[54],H2[38]} , {Pr2[21],Pr2[5],Pr2[53]} ,H3[22] ) ;
    _4G3P_G4 _4G3P_G4_87( {H2[23],H2[7],H2[55],H2[39]} , {Pr2[22],Pr2[6],Pr2[54]} ,H3[23] ) ;
    _4G3P_G4 _4G3P_G4_88( {H2[24],H2[8],H2[56],H2[40]} , {Pr2[23],Pr2[7],Pr2[55]} ,H3[24] ) ;
    _4G3P_G4 _4G3P_G4_89( {H2[25],H2[9],H2[57],H2[41]} , {Pr2[24],Pr2[8],Pr2[56]} ,H3[25] ) ;
    _4G3P_G4 _4G3P_G4_90( {H2[26],H2[10],H2[58],H2[42]} , {Pr2[25],Pr2[9],Pr2[57]} ,H3[26] ) ;
    _4G3P_G4 _4G3P_G4_91( {H2[27],H2[11],H2[59],H2[43]} , {Pr2[26],Pr2[10],Pr2[58]} ,H3[27] ) ;
    _4G3P_G4 _4G3P_G4_92( {H2[28],H2[12],H2[60],H2[44]} , {Pr2[27],Pr2[11],Pr2[59]} ,H3[28] ) ;
    _4G3P_G4 _4G3P_G4_93( {H2[29],H2[13],H2[61],H2[45]} , {Pr2[28],Pr2[12],Pr2[60]} ,H3[29] ) ;
    _4G3P_G4 _4G3P_G4_94( {H2[30],H2[14],H2[62],H2[46]} , {Pr2[29],Pr2[13],Pr2[61]} ,H3[30] ) ;
    _4G3P_G4 _4G3P_G4_95( {H2[31],H2[15],H2[63],H2[47]} , {Pr2[30],Pr2[14],Pr2[62]} ,H3[31] ) ;
    _4G3P_G4 _4G3P_G4_96( {H2[32],H2[16],H2[0],H2[48]} , {Pr2[31],Pr2[15],Pr2[63]} ,H3[32] ) ;
    _4G3P_G4 _4G3P_G4_97( {H2[33],H2[17],H2[1],H2[49]} , {Pr2[32],Pr2[16],Pr2[0]} ,H3[33] ) ;
    _4G3P_G4 _4G3P_G4_98( {H2[34],H2[18],H2[2],H2[50]} , {Pr2[33],Pr2[17],Pr2[1]} ,H3[34] ) ;
    _4G3P_G4 _4G3P_G4_99( {H2[35],H2[19],H2[3],H2[51]} , {Pr2[34],Pr2[18],Pr2[2]} ,H3[35] ) ;
    _4G3P_G4 _4G3P_G4_100( {H2[36],H2[20],H2[4],H2[52]} , {Pr2[35],Pr2[19],Pr2[3]} ,H3[36] ) ;
    _4G3P_G4 _4G3P_G4_101( {H2[37],H2[21],H2[5],H2[53]} , {Pr2[36],Pr2[20],Pr2[4]} ,H3[37] ) ;
    _4G3P_G4 _4G3P_G4_102( {H2[38],H2[22],H2[6],H2[54]} , {Pr2[37],Pr2[21],Pr2[5]} ,H3[38] ) ;
    _4G3P_G4 _4G3P_G4_103( {H2[39],H2[23],H2[7],H2[55]} , {Pr2[38],Pr2[22],Pr2[6]} ,H3[39] ) ;
    _4G3P_G4 _4G3P_G4_104( {H2[40],H2[24],H2[8],H2[56]} , {Pr2[39],Pr2[23],Pr2[7]} ,H3[40] ) ;
    _4G3P_G4 _4G3P_G4_105( {H2[41],H2[25],H2[9],H2[57]} , {Pr2[40],Pr2[24],Pr2[8]} ,H3[41] ) ;
    _4G3P_G4 _4G3P_G4_106( {H2[42],H2[26],H2[10],H2[58]} , {Pr2[41],Pr2[25],Pr2[9]} ,H3[42] ) ;
    _4G3P_G4 _4G3P_G4_107( {H2[43],H2[27],H2[11],H2[59]} , {Pr2[42],Pr2[26],Pr2[10]} ,H3[43] ) ;
    _4G3P_G4 _4G3P_G4_108( {H2[44],H2[28],H2[12],H2[60]} , {Pr2[43],Pr2[27],Pr2[11]} ,H3[44] ) ;
    _4G3P_G4 _4G3P_G4_109( {H2[45],H2[29],H2[13],H2[61]} , {Pr2[44],Pr2[28],Pr2[12]} ,H3[45] ) ;
    _4G3P_G4 _4G3P_G4_110( {H2[46],H2[30],H2[14],H2[62]} , {Pr2[45],Pr2[29],Pr2[13]} ,H3[46] ) ;
    _4G3P_G4 _4G3P_G4_111( {H2[47],H2[31],H2[15],H2[63]} , {Pr2[46],Pr2[30],Pr2[14]} ,H3[47] ) ;
    _4G3P_G4 _4G3P_G4_112( {H2[48],H2[32],H2[16],H2[0]} , {Pr2[47],Pr2[31],Pr2[15]} ,H3[48] ) ;
    _4G3P_G4 _4G3P_G4_113( {H2[49],H2[33],H2[17],H2[1]} , {Pr2[48],Pr2[32],Pr2[16]} ,H3[49] ) ;
    _4G3P_G4 _4G3P_G4_114( {H2[50],H2[34],H2[18],H2[2]} , {Pr2[49],Pr2[33],Pr2[17]} ,H3[50] ) ;
    _4G3P_G4 _4G3P_G4_115( {H2[51],H2[35],H2[19],H2[3]} , {Pr2[50],Pr2[34],Pr2[18]} ,H3[51] ) ;
    _4G3P_G4 _4G3P_G4_116( {H2[52],H2[36],H2[20],H2[4]} , {Pr2[51],Pr2[35],Pr2[19]} ,H3[52] ) ;
    _4G3P_G4 _4G3P_G4_117( {H2[53],H2[37],H2[21],H2[5]} , {Pr2[52],Pr2[36],Pr2[20]} ,H3[53] ) ;
    _4G3P_G4 _4G3P_G4_118( {H2[54],H2[38],H2[22],H2[6]} , {Pr2[53],Pr2[37],Pr2[21]} ,H3[54] ) ;
    _4G3P_G4 _4G3P_G4_119( {H2[55],H2[39],H2[23],H2[7]} , {Pr2[54],Pr2[38],Pr2[22]} ,H3[55] ) ;
    _4G3P_G4 _4G3P_G4_120( {H2[56],H2[40],H2[24],H2[8]} , {Pr2[55],Pr2[39],Pr2[23]} ,H3[56] ) ;
    _4G3P_G4 _4G3P_G4_121( {H2[57],H2[41],H2[25],H2[9]} , {Pr2[56],Pr2[40],Pr2[24]} ,H3[57] ) ;
    _4G3P_G4 _4G3P_G4_122( {H2[58],H2[42],H2[26],H2[10]} , {Pr2[57],Pr2[41],Pr2[25]} ,H3[58] ) ;
    _4G3P_G4 _4G3P_G4_123( {H2[59],H2[43],H2[27],H2[11]} , {Pr2[58],Pr2[42],Pr2[26]} ,H3[59] ) ;
    _4G3P_G4 _4G3P_G4_124( {H2[60],H2[44],H2[28],H2[12]} , {Pr2[59],Pr2[43],Pr2[27]} ,H3[60] ) ;
    _4G3P_G4 _4G3P_G4_125( {H2[61],H2[45],H2[29],H2[13]} , {Pr2[60],Pr2[44],Pr2[28]} ,H3[61] ) ;
    _4G3P_G4 _4G3P_G4_126( {H2[62],H2[46],H2[30],H2[14]} , {Pr2[61],Pr2[45],Pr2[29]} ,H3[62] ) ;
    _4G3P_G4 _4G3P_G4_127( {H2[63],H2[47],H2[31],H2[15]} , {Pr2[62],Pr2[46],Pr2[30]} ,H3[63] ) ;

    _Lsum _Lsum_0( p[63] , x[0] , H3[63] , sum[0]  ) ;
    _Lsum _Lsum_1( p[0] , x[1] , H3[0] , sum[1]  ) ;
    _Lsum _Lsum_2( p[1] , x[2] , H3[1] , sum[2]  ) ;
    _Lsum _Lsum_3( p[2] , x[3] , H3[2] , sum[3]  ) ;
    _Lsum _Lsum_4( p[3] , x[4] , H3[3] , sum[4]  ) ;
    _Lsum _Lsum_5( p[4] , x[5] , H3[4] , sum[5]  ) ;
    _Lsum _Lsum_6( p[5] , x[6] , H3[5] , sum[6]  ) ;
    _Lsum _Lsum_7( p[6] , x[7] , H3[6] , sum[7]  ) ;
    _Lsum _Lsum_8( p[7] , x[8] , H3[7] , sum[8]  ) ;
    _Lsum _Lsum_9( p[8] , x[9] , H3[8] , sum[9]  ) ;
    _Lsum _Lsum_10( p[9] , x[10] , H3[9] , sum[10]  ) ;
    _Lsum _Lsum_11( p[10] , x[11] , H3[10] , sum[11]  ) ;
    _Lsum _Lsum_12( p[11] , x[12] , H3[11] , sum[12]  ) ;
    _Lsum _Lsum_13( p[12] , x[13] , H3[12] , sum[13]  ) ;
    _Lsum _Lsum_14( p[13] , x[14] , H3[13] , sum[14]  ) ;
    _Lsum _Lsum_15( p[14] , x[15] , H3[14] , sum[15]  ) ;
    _Lsum _Lsum_16( p[15] , x[16] , H3[15] , sum[16]  ) ;
    _Lsum _Lsum_17( p[16] , x[17] , H3[16] , sum[17]  ) ;
    _Lsum _Lsum_18( p[17] , x[18] , H3[17] , sum[18]  ) ;
    _Lsum _Lsum_19( p[18] , x[19] , H3[18] , sum[19]  ) ;
    _Lsum _Lsum_20( p[19] , x[20] , H3[19] , sum[20]  ) ;
    _Lsum _Lsum_21( p[20] , x[21] , H3[20] , sum[21]  ) ;
    _Lsum _Lsum_22( p[21] , x[22] , H3[21] , sum[22]  ) ;
    _Lsum _Lsum_23( p[22] , x[23] , H3[22] , sum[23]  ) ;
    _Lsum _Lsum_24( p[23] , x[24] , H3[23] , sum[24]  ) ;
    _Lsum _Lsum_25( p[24] , x[25] , H3[24] , sum[25]  ) ;
    _Lsum _Lsum_26( p[25] , x[26] , H3[25] , sum[26]  ) ;
    _Lsum _Lsum_27( p[26] , x[27] , H3[26] , sum[27]  ) ;
    _Lsum _Lsum_28( p[27] , x[28] , H3[27] , sum[28]  ) ;
    _Lsum _Lsum_29( p[28] , x[29] , H3[28] , sum[29]  ) ;
    _Lsum _Lsum_30( p[29] , x[30] , H3[29] , sum[30]  ) ;
    _Lsum _Lsum_31( p[30] , x[31] , H3[30] , sum[31]  ) ;
    _Lsum _Lsum_32( p[31] , x[32] , H3[31] , sum[32]  ) ;
    _Lsum _Lsum_33( p[32] , x[33] , H3[32] , sum[33]  ) ;
    _Lsum _Lsum_34( p[33] , x[34] , H3[33] , sum[34]  ) ;
    _Lsum _Lsum_35( p[34] , x[35] , H3[34] , sum[35]  ) ;
    _Lsum _Lsum_36( p[35] , x[36] , H3[35] , sum[36]  ) ;
    _Lsum _Lsum_37( p[36] , x[37] , H3[36] , sum[37]  ) ;
    _Lsum _Lsum_38( p[37] , x[38] , H3[37] , sum[38]  ) ;
    _Lsum _Lsum_39( p[38] , x[39] , H3[38] , sum[39]  ) ;
    _Lsum _Lsum_40( p[39] , x[40] , H3[39] , sum[40]  ) ;
    _Lsum _Lsum_41( p[40] , x[41] , H3[40] , sum[41]  ) ;
    _Lsum _Lsum_42( p[41] , x[42] , H3[41] , sum[42]  ) ;
    _Lsum _Lsum_43( p[42] , x[43] , H3[42] , sum[43]  ) ;
    _Lsum _Lsum_44( p[43] , x[44] , H3[43] , sum[44]  ) ;
    _Lsum _Lsum_45( p[44] , x[45] , H3[44] , sum[45]  ) ;
    _Lsum _Lsum_46( p[45] , x[46] , H3[45] , sum[46]  ) ;
    _Lsum _Lsum_47( p[46] , x[47] , H3[46] , sum[47]  ) ;
    _Lsum _Lsum_48( p[47] , x[48] , H3[47] , sum[48]  ) ;
    _Lsum _Lsum_49( p[48] , x[49] , H3[48] , sum[49]  ) ;
    _Lsum _Lsum_50( p[49] , x[50] , H3[49] , sum[50]  ) ;
    _Lsum _Lsum_51( p[50] , x[51] , H3[50] , sum[51]  ) ;
    _Lsum _Lsum_52( p[51] , x[52] , H3[51] , sum[52]  ) ;
    _Lsum _Lsum_53( p[52] , x[53] , H3[52] , sum[53]  ) ;
    _Lsum _Lsum_54( p[53] , x[54] , H3[53] , sum[54]  ) ;
    _Lsum _Lsum_55( p[54] , x[55] , H3[54] , sum[55]  ) ;
    _Lsum _Lsum_56( p[55] , x[56] , H3[55] , sum[56]  ) ;
    _Lsum _Lsum_57( p[56] , x[57] , H3[56] , sum[57]  ) ;
    _Lsum _Lsum_58( p[57] , x[58] , H3[57] , sum[58]  ) ;
    _Lsum _Lsum_59( p[58] , x[59] , H3[58] , sum[59]  ) ;
    _Lsum _Lsum_60( p[59] , x[60] , H3[59] , sum[60]  ) ;
    _Lsum _Lsum_61( p[60] , x[61] , H3[60] , sum[61]  ) ;
    _Lsum _Lsum_62( p[61] , x[62] , H3[61] , sum[62]  ) ;
    _Lsum _Lsum_63( p[62] , x[63] , H3[62] , sum[63]  ) ;

endmodule
