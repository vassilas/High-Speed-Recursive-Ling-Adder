module J8_node_adder(a, b, sum);
    input [7:0]a;
    input [7:0]b;
    output [7:0]sum;
    wire [7:0]g ;
    wire [7:0]p ;
    wire [7:0]x ;
    wire [7:0]R1 ;
    wire [7:0]R2 ;
    wire [7:0]Q1 ;
    wire [7:0]D1 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;

    _2g_R2 _2g_R2_0( {g[0],g[7] } , R1[0] ) ;
    _2g_R2 _2g_R2_1( {g[1],g[0] } , R1[1] ) ;
    _2g_R2 _2g_R2_2( {g[2],g[1] } , R1[2] ) ;
    _2g_R2 _2g_R2_3( {g[3],g[2] } , R1[3] ) ;
    _2g_R2 _2g_R2_4( {g[4],g[3] } , R1[4] ) ;
    _2g_R2 _2g_R2_5( {g[5],g[4] } , R1[5] ) ;
    _2g_R2 _2g_R2_6( {g[6],g[5] } , R1[6] ) ;
    _2g_R2 _2g_R2_7( {g[7],g[6] } , R1[7] ) ;

    _2p_Q2 _2p_Q2_0( {p[0],p[7] } , Q1[0] ) ;
    _2p_Q2 _2p_Q2_1( {p[1],p[0] } , Q1[1] ) ;
    _2p_Q2 _2p_Q2_2( {p[2],p[1] } , Q1[2] ) ;
    _2p_Q2 _2p_Q2_3( {p[3],p[2] } , Q1[3] ) ;
    _2p_Q2 _2p_Q2_4( {p[4],p[3] } , Q1[4] ) ;
    _2p_Q2 _2p_Q2_5( {p[5],p[4] } , Q1[5] ) ;
    _2p_Q2 _2p_Q2_6( {p[6],p[5] } , Q1[6] ) ;
    _2p_Q2 _2p_Q2_7( {p[7],p[6] } , Q1[7] ) ;

    _4R2Q_R4 _4R2Q_R4_0( {R1[0],R1[6],R1[4],R1[2] }, {Q1[5],Q1[3]} ,R2[0] ) ;
    _4R2Q_R4 _4R2Q_R4_1( {R1[1],R1[7],R1[5],R1[3] }, {Q1[6],Q1[4]} ,R2[1] ) ;
    _4R2Q_R4 _4R2Q_R4_2( {R1[2],R1[0],R1[6],R1[4] }, {Q1[7],Q1[5]} ,R2[2] ) ;
    _4R2Q_R4 _4R2Q_R4_3( {R1[3],R1[1],R1[7],R1[5] }, {Q1[0],Q1[6]} ,R2[3] ) ;
    _4R2Q_R4 _4R2Q_R4_4( {R1[4],R1[2],R1[0],R1[6] }, {Q1[1],Q1[7]} ,R2[4] ) ;
    _4R2Q_R4 _4R2Q_R4_5( {R1[5],R1[3],R1[1],R1[7] }, {Q1[2],Q1[0]} ,R2[5] ) ;
    _4R2Q_R4 _4R2Q_R4_6( {R1[6],R1[4],R1[2],R1[0] }, {Q1[3],Q1[1]} ,R2[6] ) ;
    _4R2Q_R4 _4R2Q_R4_7( {R1[7],R1[5],R1[3],R1[1] }, {Q1[4],Q1[2]} ,R2[7] ) ;

    _D64_1 _D64_1_0( {p[0],p[7],p[6]}, {g[0],g[7]}, D1[0] ) ;
    _D64_1 _D64_1_1( {p[1],p[0],p[7]}, {g[1],g[0]}, D1[1] ) ;
    _D64_1 _D64_1_2( {p[2],p[1],p[0]}, {g[2],g[1]}, D1[2] ) ;
    _D64_1 _D64_1_3( {p[3],p[2],p[1]}, {g[3],g[2]}, D1[3] ) ;
    _D64_1 _D64_1_4( {p[4],p[3],p[2]}, {g[4],g[3]}, D1[4] ) ;
    _D64_1 _D64_1_5( {p[5],p[4],p[3]}, {g[5],g[4]}, D1[5] ) ;
    _D64_1 _D64_1_6( {p[6],p[5],p[4]}, {g[6],g[5]}, D1[6] ) ;
    _D64_1 _D64_1_7( {p[7],p[6],p[5]}, {g[7],g[6]}, D1[7] ) ;

    _Jsum _Jsum_0( R2[7], D1[7] , x[0] , sum[0] ) ;
    _Jsum _Jsum_1( R2[0], D1[0] , x[1] , sum[1] ) ;
    _Jsum _Jsum_2( R2[1], D1[1] , x[2] , sum[2] ) ;
    _Jsum _Jsum_3( R2[2], D1[2] , x[3] , sum[3] ) ;
    _Jsum _Jsum_4( R2[3], D1[3] , x[4] , sum[4] ) ;
    _Jsum _Jsum_5( R2[4], D1[4] , x[5] , sum[5] ) ;
    _Jsum _Jsum_6( R2[5], D1[5] , x[6] , sum[6] ) ;
    _Jsum _Jsum_7( R2[6], D1[6] , x[7] , sum[7] ) ;

endmodule
