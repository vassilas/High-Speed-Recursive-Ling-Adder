module L16_node_adder(a, b, sum);
    input [15:0]a;
    input [15:0]b;
    output [15:0]sum;
    wire [15:0]g ;
    wire [15:0]p ;
    wire [15:0]x ;
    wire [15:0]H1 ;
    wire [15:0]H2 ;
    wire [15:0]Pr1 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;

    _4g2p_H4 _4g2p_H4_0( {g[0],g[15],g[14],g[13]} ,{p[15],p[14]} , H1[0] ) ;
    _4g2p_H4 _4g2p_H4_1( {g[1],g[0],g[15],g[14]} ,{p[0],p[15]} , H1[1] ) ;
    _4g2p_H4 _4g2p_H4_2( {g[2],g[1],g[0],g[15]} ,{p[1],p[0]} , H1[2] ) ;
    _4g2p_H4 _4g2p_H4_3( {g[3],g[2],g[1],g[0]} ,{p[2],p[1]} , H1[3] ) ;
    _4g2p_H4 _4g2p_H4_4( {g[4],g[3],g[2],g[1]} ,{p[3],p[2]} , H1[4] ) ;
    _4g2p_H4 _4g2p_H4_5( {g[5],g[4],g[3],g[2]} ,{p[4],p[3]} , H1[5] ) ;
    _4g2p_H4 _4g2p_H4_6( {g[6],g[5],g[4],g[3]} ,{p[5],p[4]} , H1[6] ) ;
    _4g2p_H4 _4g2p_H4_7( {g[7],g[6],g[5],g[4]} ,{p[6],p[5]} , H1[7] ) ;
    _4g2p_H4 _4g2p_H4_8( {g[8],g[7],g[6],g[5]} ,{p[7],p[6]} , H1[8] ) ;
    _4g2p_H4 _4g2p_H4_9( {g[9],g[8],g[7],g[6]} ,{p[8],p[7]} , H1[9] ) ;
    _4g2p_H4 _4g2p_H4_10( {g[10],g[9],g[8],g[7]} ,{p[9],p[8]} , H1[10] ) ;
    _4g2p_H4 _4g2p_H4_11( {g[11],g[10],g[9],g[8]} ,{p[10],p[9]} , H1[11] ) ;
    _4g2p_H4 _4g2p_H4_12( {g[12],g[11],g[10],g[9]} ,{p[11],p[10]} , H1[12] ) ;
    _4g2p_H4 _4g2p_H4_13( {g[13],g[12],g[11],g[10]} ,{p[12],p[11]} , H1[13] ) ;
    _4g2p_H4 _4g2p_H4_14( {g[14],g[13],g[12],g[11]} ,{p[13],p[12]} , H1[14] ) ;
    _4g2p_H4 _4g2p_H4_15( {g[15],g[14],g[13],g[12]} ,{p[14],p[13]} , H1[15] ) ;

    _P4 _P4_0( {p[0],p[15],p[14],p[13]} ,Pr1[0] ) ;
    _P4 _P4_1( {p[1],p[0],p[15],p[14]} ,Pr1[1] ) ;
    _P4 _P4_2( {p[2],p[1],p[0],p[15]} ,Pr1[2] ) ;
    _P4 _P4_3( {p[3],p[2],p[1],p[0]} ,Pr1[3] ) ;
    _P4 _P4_4( {p[4],p[3],p[2],p[1]} ,Pr1[4] ) ;
    _P4 _P4_5( {p[5],p[4],p[3],p[2]} ,Pr1[5] ) ;
    _P4 _P4_6( {p[6],p[5],p[4],p[3]} ,Pr1[6] ) ;
    _P4 _P4_7( {p[7],p[6],p[5],p[4]} ,Pr1[7] ) ;
    _P4 _P4_8( {p[8],p[7],p[6],p[5]} ,Pr1[8] ) ;
    _P4 _P4_9( {p[9],p[8],p[7],p[6]} ,Pr1[9] ) ;
    _P4 _P4_10( {p[10],p[9],p[8],p[7]} ,Pr1[10] ) ;
    _P4 _P4_11( {p[11],p[10],p[9],p[8]} ,Pr1[11] ) ;
    _P4 _P4_12( {p[12],p[11],p[10],p[9]} ,Pr1[12] ) ;
    _P4 _P4_13( {p[13],p[12],p[11],p[10]} ,Pr1[13] ) ;
    _P4 _P4_14( {p[14],p[13],p[12],p[11]} ,Pr1[14] ) ;
    _P4 _P4_15( {p[15],p[14],p[13],p[12]} ,Pr1[15] ) ;

    _4G3P_G4 _4G3P_G4_0( {H1[0],H1[12],H1[8],H1[4]} , {Pr1[15],Pr1[11],Pr1[7]} ,H2[0] ) ;
    _4G3P_G4 _4G3P_G4_1( {H1[1],H1[13],H1[9],H1[5]} , {Pr1[0],Pr1[12],Pr1[8]} ,H2[1] ) ;
    _4G3P_G4 _4G3P_G4_2( {H1[2],H1[14],H1[10],H1[6]} , {Pr1[1],Pr1[13],Pr1[9]} ,H2[2] ) ;
    _4G3P_G4 _4G3P_G4_3( {H1[3],H1[15],H1[11],H1[7]} , {Pr1[2],Pr1[14],Pr1[10]} ,H2[3] ) ;
    _4G3P_G4 _4G3P_G4_4( {H1[4],H1[0],H1[12],H1[8]} , {Pr1[3],Pr1[15],Pr1[11]} ,H2[4] ) ;
    _4G3P_G4 _4G3P_G4_5( {H1[5],H1[1],H1[13],H1[9]} , {Pr1[4],Pr1[0],Pr1[12]} ,H2[5] ) ;
    _4G3P_G4 _4G3P_G4_6( {H1[6],H1[2],H1[14],H1[10]} , {Pr1[5],Pr1[1],Pr1[13]} ,H2[6] ) ;
    _4G3P_G4 _4G3P_G4_7( {H1[7],H1[3],H1[15],H1[11]} , {Pr1[6],Pr1[2],Pr1[14]} ,H2[7] ) ;
    _4G3P_G4 _4G3P_G4_8( {H1[8],H1[4],H1[0],H1[12]} , {Pr1[7],Pr1[3],Pr1[15]} ,H2[8] ) ;
    _4G3P_G4 _4G3P_G4_9( {H1[9],H1[5],H1[1],H1[13]} , {Pr1[8],Pr1[4],Pr1[0]} ,H2[9] ) ;
    _4G3P_G4 _4G3P_G4_10( {H1[10],H1[6],H1[2],H1[14]} , {Pr1[9],Pr1[5],Pr1[1]} ,H2[10] ) ;
    _4G3P_G4 _4G3P_G4_11( {H1[11],H1[7],H1[3],H1[15]} , {Pr1[10],Pr1[6],Pr1[2]} ,H2[11] ) ;
    _4G3P_G4 _4G3P_G4_12( {H1[12],H1[8],H1[4],H1[0]} , {Pr1[11],Pr1[7],Pr1[3]} ,H2[12] ) ;
    _4G3P_G4 _4G3P_G4_13( {H1[13],H1[9],H1[5],H1[1]} , {Pr1[12],Pr1[8],Pr1[4]} ,H2[13] ) ;
    _4G3P_G4 _4G3P_G4_14( {H1[14],H1[10],H1[6],H1[2]} , {Pr1[13],Pr1[9],Pr1[5]} ,H2[14] ) ;
    _4G3P_G4 _4G3P_G4_15( {H1[15],H1[11],H1[7],H1[3]} , {Pr1[14],Pr1[10],Pr1[6]} ,H2[15] ) ;

    _Lsum _Lsum_0( p[15] , x[0] , H2[15] , sum[0]  ) ;
    _Lsum _Lsum_1( p[0] , x[1] , H2[0] , sum[1]  ) ;
    _Lsum _Lsum_2( p[1] , x[2] , H2[1] , sum[2]  ) ;
    _Lsum _Lsum_3( p[2] , x[3] , H2[2] , sum[3]  ) ;
    _Lsum _Lsum_4( p[3] , x[4] , H2[3] , sum[4]  ) ;
    _Lsum _Lsum_5( p[4] , x[5] , H2[4] , sum[5]  ) ;
    _Lsum _Lsum_6( p[5] , x[6] , H2[5] , sum[6]  ) ;
    _Lsum _Lsum_7( p[6] , x[7] , H2[6] , sum[7]  ) ;
    _Lsum _Lsum_8( p[7] , x[8] , H2[7] , sum[8]  ) ;
    _Lsum _Lsum_9( p[8] , x[9] , H2[8] , sum[9]  ) ;
    _Lsum _Lsum_10( p[9] , x[10] , H2[9] , sum[10]  ) ;
    _Lsum _Lsum_11( p[10] , x[11] , H2[10] , sum[11]  ) ;
    _Lsum _Lsum_12( p[11] , x[12] , H2[11] , sum[12]  ) ;
    _Lsum _Lsum_13( p[12] , x[13] , H2[12] , sum[13]  ) ;
    _Lsum _Lsum_14( p[13] , x[14] , H2[13] , sum[14]  ) ;
    _Lsum _Lsum_15( p[14] , x[15] , H2[14] , sum[15]  ) ;

endmodule
