module P16_node_adder(a, b, sum);
    input [15:0]a;
    input [15:0]b;
    output [15:0]sum;
    wire [15:0]g ;
    wire [15:0]p ;
    wire [15:0]x ;
    wire [15:0]G1 ;
    wire [15:0]G2 ;
    wire [15:0]Pr1 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;

    _4G3P_G4 _4G3P_G4_3( {g[3],g[2],g[1],g[0]} , {p[3],p[2],p[1]} ,G1[3] ) ;
    _4G3P_G4 _4G3P_G4_7( {g[7],g[6],g[5],g[4]} , {p[7],p[6],p[5]} ,G1[7] ) ;
    _4G3P_G4 _4G3P_G4_11( {g[11],g[10],g[9],g[8]} , {p[11],p[10],p[9]} ,G1[11] ) ;
    _4G3P_G4 _4G3P_G4_15( {g[15],g[14],g[13],g[12]} , {p[15],p[14],p[13]} ,G1[15] ) ;

    _P4 _P4_3( {p[3],p[2],p[1],p[0]} ,Pr1[3] ) ;
    _P4 _P4_7( {p[7],p[6],p[5],p[4]} ,Pr1[7] ) ;
    _P4 _P4_11( {p[11],p[10],p[9],p[8]} ,Pr1[11] ) ;
    _P4 _P4_15( {p[15],p[14],p[13],p[12]} ,Pr1[15] ) ;

    _4G3P_G4 _4G3P_G4_19( {G1[3],G1[15],G1[11],G1[7]} , {Pr1[3],Pr1[15],Pr1[11]} ,G2[3] ) ;
    _4G3P_G4 _4G3P_G4_23( {G1[7],G1[3],G1[15],G1[11]} , {Pr1[7],Pr1[3],Pr1[15]} ,G2[7] ) ;
    _4G3P_G4 _4G3P_G4_27( {G1[11],G1[7],G1[3],G1[15]} , {Pr1[11],Pr1[7],Pr1[3]} ,G2[11] ) ;
    _4G3P_G4 _4G3P_G4_31( {G1[15],G1[11],G1[7],G1[3]} , {Pr1[15],Pr1[11],Pr1[7]} ,G2[15] ) ;

    _Psum_sparse4 _Psum_sparse4_0( {x[3],x[2],x[1],x[0]} ,  {g[2],g[1],g[0]} , {p[2],p[1],p[0]} , G2[15] , {sum[3],sum[2],sum[1],sum[0]} ) ;
    _Psum_sparse4 _Psum_sparse4_4( {x[7],x[6],x[5],x[4]} ,  {g[6],g[5],g[4]} , {p[6],p[5],p[4]} , G2[3] , {sum[7],sum[6],sum[5],sum[4]} ) ;
    _Psum_sparse4 _Psum_sparse4_8( {x[11],x[10],x[9],x[8]} ,  {g[10],g[9],g[8]} , {p[10],p[9],p[8]} , G2[7] , {sum[11],sum[10],sum[9],sum[8]} ) ;
    _Psum_sparse4 _Psum_sparse4_12( {x[15],x[14],x[13],x[12]} ,  {g[14],g[13],g[12]} , {p[14],p[13],p[12]} , G2[11] , {sum[15],sum[14],sum[13],sum[12]} ) ;

endmodule
