module P64_node_adder(a, b, sum);
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    wire [63:0]g ;
    wire [63:0]p ;
    wire [63:0]x ;
    wire [63:0]G1 ;
    wire [63:0]G2 ;
    wire [63:0]G3 ;
    wire [63:0]Pr1 ;
    wire [63:0]Pr2 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;
    _gpx _gpx_16	(a[16],	b[16],	g[16], 	p[16], 	x[16]) ;
    _gpx _gpx_17	(a[17],	b[17],	g[17], 	p[17], 	x[17]) ;
    _gpx _gpx_18	(a[18],	b[18],	g[18], 	p[18], 	x[18]) ;
    _gpx _gpx_19	(a[19],	b[19],	g[19], 	p[19], 	x[19]) ;
    _gpx _gpx_20	(a[20],	b[20],	g[20], 	p[20], 	x[20]) ;
    _gpx _gpx_21	(a[21],	b[21],	g[21], 	p[21], 	x[21]) ;
    _gpx _gpx_22	(a[22],	b[22],	g[22], 	p[22], 	x[22]) ;
    _gpx _gpx_23	(a[23],	b[23],	g[23], 	p[23], 	x[23]) ;
    _gpx _gpx_24	(a[24],	b[24],	g[24], 	p[24], 	x[24]) ;
    _gpx _gpx_25	(a[25],	b[25],	g[25], 	p[25], 	x[25]) ;
    _gpx _gpx_26	(a[26],	b[26],	g[26], 	p[26], 	x[26]) ;
    _gpx _gpx_27	(a[27],	b[27],	g[27], 	p[27], 	x[27]) ;
    _gpx _gpx_28	(a[28],	b[28],	g[28], 	p[28], 	x[28]) ;
    _gpx _gpx_29	(a[29],	b[29],	g[29], 	p[29], 	x[29]) ;
    _gpx _gpx_30	(a[30],	b[30],	g[30], 	p[30], 	x[30]) ;
    _gpx _gpx_31	(a[31],	b[31],	g[31], 	p[31], 	x[31]) ;
    _gpx _gpx_32	(a[32],	b[32],	g[32], 	p[32], 	x[32]) ;
    _gpx _gpx_33	(a[33],	b[33],	g[33], 	p[33], 	x[33]) ;
    _gpx _gpx_34	(a[34],	b[34],	g[34], 	p[34], 	x[34]) ;
    _gpx _gpx_35	(a[35],	b[35],	g[35], 	p[35], 	x[35]) ;
    _gpx _gpx_36	(a[36],	b[36],	g[36], 	p[36], 	x[36]) ;
    _gpx _gpx_37	(a[37],	b[37],	g[37], 	p[37], 	x[37]) ;
    _gpx _gpx_38	(a[38],	b[38],	g[38], 	p[38], 	x[38]) ;
    _gpx _gpx_39	(a[39],	b[39],	g[39], 	p[39], 	x[39]) ;
    _gpx _gpx_40	(a[40],	b[40],	g[40], 	p[40], 	x[40]) ;
    _gpx _gpx_41	(a[41],	b[41],	g[41], 	p[41], 	x[41]) ;
    _gpx _gpx_42	(a[42],	b[42],	g[42], 	p[42], 	x[42]) ;
    _gpx _gpx_43	(a[43],	b[43],	g[43], 	p[43], 	x[43]) ;
    _gpx _gpx_44	(a[44],	b[44],	g[44], 	p[44], 	x[44]) ;
    _gpx _gpx_45	(a[45],	b[45],	g[45], 	p[45], 	x[45]) ;
    _gpx _gpx_46	(a[46],	b[46],	g[46], 	p[46], 	x[46]) ;
    _gpx _gpx_47	(a[47],	b[47],	g[47], 	p[47], 	x[47]) ;
    _gpx _gpx_48	(a[48],	b[48],	g[48], 	p[48], 	x[48]) ;
    _gpx _gpx_49	(a[49],	b[49],	g[49], 	p[49], 	x[49]) ;
    _gpx _gpx_50	(a[50],	b[50],	g[50], 	p[50], 	x[50]) ;
    _gpx _gpx_51	(a[51],	b[51],	g[51], 	p[51], 	x[51]) ;
    _gpx _gpx_52	(a[52],	b[52],	g[52], 	p[52], 	x[52]) ;
    _gpx _gpx_53	(a[53],	b[53],	g[53], 	p[53], 	x[53]) ;
    _gpx _gpx_54	(a[54],	b[54],	g[54], 	p[54], 	x[54]) ;
    _gpx _gpx_55	(a[55],	b[55],	g[55], 	p[55], 	x[55]) ;
    _gpx _gpx_56	(a[56],	b[56],	g[56], 	p[56], 	x[56]) ;
    _gpx _gpx_57	(a[57],	b[57],	g[57], 	p[57], 	x[57]) ;
    _gpx _gpx_58	(a[58],	b[58],	g[58], 	p[58], 	x[58]) ;
    _gpx _gpx_59	(a[59],	b[59],	g[59], 	p[59], 	x[59]) ;
    _gpx _gpx_60	(a[60],	b[60],	g[60], 	p[60], 	x[60]) ;
    _gpx _gpx_61	(a[61],	b[61],	g[61], 	p[61], 	x[61]) ;
    _gpx _gpx_62	(a[62],	b[62],	g[62], 	p[62], 	x[62]) ;
    _gpx _gpx_63	(a[63],	b[63],	g[63], 	p[63], 	x[63]) ;

    _4G3P_G4 _4G3P_G4_3( {g[3],g[2],g[1],g[0]} , {p[3],p[2],p[1]} ,G1[3] ) ;
    _4G3P_G4 _4G3P_G4_7( {g[7],g[6],g[5],g[4]} , {p[7],p[6],p[5]} ,G1[7] ) ;
    _4G3P_G4 _4G3P_G4_11( {g[11],g[10],g[9],g[8]} , {p[11],p[10],p[9]} ,G1[11] ) ;
    _4G3P_G4 _4G3P_G4_15( {g[15],g[14],g[13],g[12]} , {p[15],p[14],p[13]} ,G1[15] ) ;
    _4G3P_G4 _4G3P_G4_19( {g[19],g[18],g[17],g[16]} , {p[19],p[18],p[17]} ,G1[19] ) ;
    _4G3P_G4 _4G3P_G4_23( {g[23],g[22],g[21],g[20]} , {p[23],p[22],p[21]} ,G1[23] ) ;
    _4G3P_G4 _4G3P_G4_27( {g[27],g[26],g[25],g[24]} , {p[27],p[26],p[25]} ,G1[27] ) ;
    _4G3P_G4 _4G3P_G4_31( {g[31],g[30],g[29],g[28]} , {p[31],p[30],p[29]} ,G1[31] ) ;
    _4G3P_G4 _4G3P_G4_35( {g[35],g[34],g[33],g[32]} , {p[35],p[34],p[33]} ,G1[35] ) ;
    _4G3P_G4 _4G3P_G4_39( {g[39],g[38],g[37],g[36]} , {p[39],p[38],p[37]} ,G1[39] ) ;
    _4G3P_G4 _4G3P_G4_43( {g[43],g[42],g[41],g[40]} , {p[43],p[42],p[41]} ,G1[43] ) ;
    _4G3P_G4 _4G3P_G4_47( {g[47],g[46],g[45],g[44]} , {p[47],p[46],p[45]} ,G1[47] ) ;
    _4G3P_G4 _4G3P_G4_51( {g[51],g[50],g[49],g[48]} , {p[51],p[50],p[49]} ,G1[51] ) ;
    _4G3P_G4 _4G3P_G4_55( {g[55],g[54],g[53],g[52]} , {p[55],p[54],p[53]} ,G1[55] ) ;
    _4G3P_G4 _4G3P_G4_59( {g[59],g[58],g[57],g[56]} , {p[59],p[58],p[57]} ,G1[59] ) ;
    _4G3P_G4 _4G3P_G4_63( {g[63],g[62],g[61],g[60]} , {p[63],p[62],p[61]} ,G1[63] ) ;

    _P4 _P4_3( {p[3],p[2],p[1],p[0]} ,Pr1[3] ) ;
    _P4 _P4_7( {p[7],p[6],p[5],p[4]} ,Pr1[7] ) ;
    _P4 _P4_11( {p[11],p[10],p[9],p[8]} ,Pr1[11] ) ;
    _P4 _P4_15( {p[15],p[14],p[13],p[12]} ,Pr1[15] ) ;
    _P4 _P4_19( {p[19],p[18],p[17],p[16]} ,Pr1[19] ) ;
    _P4 _P4_23( {p[23],p[22],p[21],p[20]} ,Pr1[23] ) ;
    _P4 _P4_27( {p[27],p[26],p[25],p[24]} ,Pr1[27] ) ;
    _P4 _P4_31( {p[31],p[30],p[29],p[28]} ,Pr1[31] ) ;
    _P4 _P4_35( {p[35],p[34],p[33],p[32]} ,Pr1[35] ) ;
    _P4 _P4_39( {p[39],p[38],p[37],p[36]} ,Pr1[39] ) ;
    _P4 _P4_43( {p[43],p[42],p[41],p[40]} ,Pr1[43] ) ;
    _P4 _P4_47( {p[47],p[46],p[45],p[44]} ,Pr1[47] ) ;
    _P4 _P4_51( {p[51],p[50],p[49],p[48]} ,Pr1[51] ) ;
    _P4 _P4_55( {p[55],p[54],p[53],p[52]} ,Pr1[55] ) ;
    _P4 _P4_59( {p[59],p[58],p[57],p[56]} ,Pr1[59] ) ;
    _P4 _P4_63( {p[63],p[62],p[61],p[60]} ,Pr1[63] ) ;

    _4G3P_G4 _4G3P_G4_67( {G1[3],G1[63],G1[59],G1[55]} , {Pr1[3],Pr1[63],Pr1[59]} ,G2[3] ) ;
    _4G3P_G4 _4G3P_G4_71( {G1[7],G1[3],G1[63],G1[59]} , {Pr1[7],Pr1[3],Pr1[63]} ,G2[7] ) ;
    _4G3P_G4 _4G3P_G4_75( {G1[11],G1[7],G1[3],G1[63]} , {Pr1[11],Pr1[7],Pr1[3]} ,G2[11] ) ;
    _4G3P_G4 _4G3P_G4_79( {G1[15],G1[11],G1[7],G1[3]} , {Pr1[15],Pr1[11],Pr1[7]} ,G2[15] ) ;
    _4G3P_G4 _4G3P_G4_83( {G1[19],G1[15],G1[11],G1[7]} , {Pr1[19],Pr1[15],Pr1[11]} ,G2[19] ) ;
    _4G3P_G4 _4G3P_G4_87( {G1[23],G1[19],G1[15],G1[11]} , {Pr1[23],Pr1[19],Pr1[15]} ,G2[23] ) ;
    _4G3P_G4 _4G3P_G4_91( {G1[27],G1[23],G1[19],G1[15]} , {Pr1[27],Pr1[23],Pr1[19]} ,G2[27] ) ;
    _4G3P_G4 _4G3P_G4_95( {G1[31],G1[27],G1[23],G1[19]} , {Pr1[31],Pr1[27],Pr1[23]} ,G2[31] ) ;
    _4G3P_G4 _4G3P_G4_99( {G1[35],G1[31],G1[27],G1[23]} , {Pr1[35],Pr1[31],Pr1[27]} ,G2[35] ) ;
    _4G3P_G4 _4G3P_G4_103( {G1[39],G1[35],G1[31],G1[27]} , {Pr1[39],Pr1[35],Pr1[31]} ,G2[39] ) ;
    _4G3P_G4 _4G3P_G4_107( {G1[43],G1[39],G1[35],G1[31]} , {Pr1[43],Pr1[39],Pr1[35]} ,G2[43] ) ;
    _4G3P_G4 _4G3P_G4_111( {G1[47],G1[43],G1[39],G1[35]} , {Pr1[47],Pr1[43],Pr1[39]} ,G2[47] ) ;
    _4G3P_G4 _4G3P_G4_115( {G1[51],G1[47],G1[43],G1[39]} , {Pr1[51],Pr1[47],Pr1[43]} ,G2[51] ) ;
    _4G3P_G4 _4G3P_G4_119( {G1[55],G1[51],G1[47],G1[43]} , {Pr1[55],Pr1[51],Pr1[47]} ,G2[55] ) ;
    _4G3P_G4 _4G3P_G4_123( {G1[59],G1[55],G1[51],G1[47]} , {Pr1[59],Pr1[55],Pr1[51]} ,G2[59] ) ;
    _4G3P_G4 _4G3P_G4_127( {G1[63],G1[59],G1[55],G1[51]} , {Pr1[63],Pr1[59],Pr1[55]} ,G2[63] ) ;

    _P4 _P4_67( {Pr1[3],Pr1[63],Pr1[59],Pr1[55]} ,Pr2[3] ) ;
    _P4 _P4_71( {Pr1[7],Pr1[3],Pr1[63],Pr1[59]} ,Pr2[7] ) ;
    _P4 _P4_75( {Pr1[11],Pr1[7],Pr1[3],Pr1[63]} ,Pr2[11] ) ;
    _P4 _P4_79( {Pr1[15],Pr1[11],Pr1[7],Pr1[3]} ,Pr2[15] ) ;
    _P4 _P4_83( {Pr1[19],Pr1[15],Pr1[11],Pr1[7]} ,Pr2[19] ) ;
    _P4 _P4_87( {Pr1[23],Pr1[19],Pr1[15],Pr1[11]} ,Pr2[23] ) ;
    _P4 _P4_91( {Pr1[27],Pr1[23],Pr1[19],Pr1[15]} ,Pr2[27] ) ;
    _P4 _P4_95( {Pr1[31],Pr1[27],Pr1[23],Pr1[19]} ,Pr2[31] ) ;
    _P4 _P4_99( {Pr1[35],Pr1[31],Pr1[27],Pr1[23]} ,Pr2[35] ) ;
    _P4 _P4_103( {Pr1[39],Pr1[35],Pr1[31],Pr1[27]} ,Pr2[39] ) ;
    _P4 _P4_107( {Pr1[43],Pr1[39],Pr1[35],Pr1[31]} ,Pr2[43] ) ;
    _P4 _P4_111( {Pr1[47],Pr1[43],Pr1[39],Pr1[35]} ,Pr2[47] ) ;
    _P4 _P4_115( {Pr1[51],Pr1[47],Pr1[43],Pr1[39]} ,Pr2[51] ) ;
    _P4 _P4_119( {Pr1[55],Pr1[51],Pr1[47],Pr1[43]} ,Pr2[55] ) ;
    _P4 _P4_123( {Pr1[59],Pr1[55],Pr1[51],Pr1[47]} ,Pr2[59] ) ;
    _P4 _P4_127( {Pr1[63],Pr1[59],Pr1[55],Pr1[51]} ,Pr2[63] ) ;

    _4G3P_G4 _4G3P_G4_131( {G2[3],G2[51],G2[35],G2[19]} , {Pr2[3],Pr2[51],Pr2[35]} ,G3[3] ) ;
    _4G3P_G4 _4G3P_G4_135( {G2[7],G2[55],G2[39],G2[23]} , {Pr2[7],Pr2[55],Pr2[39]} ,G3[7] ) ;
    _4G3P_G4 _4G3P_G4_139( {G2[11],G2[59],G2[43],G2[27]} , {Pr2[11],Pr2[59],Pr2[43]} ,G3[11] ) ;
    _4G3P_G4 _4G3P_G4_143( {G2[15],G2[63],G2[47],G2[31]} , {Pr2[15],Pr2[63],Pr2[47]} ,G3[15] ) ;
    _4G3P_G4 _4G3P_G4_147( {G2[19],G2[3],G2[51],G2[35]} , {Pr2[19],Pr2[3],Pr2[51]} ,G3[19] ) ;
    _4G3P_G4 _4G3P_G4_151( {G2[23],G2[7],G2[55],G2[39]} , {Pr2[23],Pr2[7],Pr2[55]} ,G3[23] ) ;
    _4G3P_G4 _4G3P_G4_155( {G2[27],G2[11],G2[59],G2[43]} , {Pr2[27],Pr2[11],Pr2[59]} ,G3[27] ) ;
    _4G3P_G4 _4G3P_G4_159( {G2[31],G2[15],G2[63],G2[47]} , {Pr2[31],Pr2[15],Pr2[63]} ,G3[31] ) ;
    _4G3P_G4 _4G3P_G4_163( {G2[35],G2[19],G2[3],G2[51]} , {Pr2[35],Pr2[19],Pr2[3]} ,G3[35] ) ;
    _4G3P_G4 _4G3P_G4_167( {G2[39],G2[23],G2[7],G2[55]} , {Pr2[39],Pr2[23],Pr2[7]} ,G3[39] ) ;
    _4G3P_G4 _4G3P_G4_171( {G2[43],G2[27],G2[11],G2[59]} , {Pr2[43],Pr2[27],Pr2[11]} ,G3[43] ) ;
    _4G3P_G4 _4G3P_G4_175( {G2[47],G2[31],G2[15],G2[63]} , {Pr2[47],Pr2[31],Pr2[15]} ,G3[47] ) ;
    _4G3P_G4 _4G3P_G4_179( {G2[51],G2[35],G2[19],G2[3]} , {Pr2[51],Pr2[35],Pr2[19]} ,G3[51] ) ;
    _4G3P_G4 _4G3P_G4_183( {G2[55],G2[39],G2[23],G2[7]} , {Pr2[55],Pr2[39],Pr2[23]} ,G3[55] ) ;
    _4G3P_G4 _4G3P_G4_187( {G2[59],G2[43],G2[27],G2[11]} , {Pr2[59],Pr2[43],Pr2[27]} ,G3[59] ) ;
    _4G3P_G4 _4G3P_G4_191( {G2[63],G2[47],G2[31],G2[15]} , {Pr2[63],Pr2[47],Pr2[31]} ,G3[63] ) ;

    _Psum_sparse4 _Psum_sparse4_0( {x[3],x[2],x[1],x[0]} ,  {g[2],g[1],g[0]} , {p[2],p[1],p[0]} , G3[63] , {sum[3],sum[2],sum[1],sum[0]} ) ;
    _Psum_sparse4 _Psum_sparse4_4( {x[7],x[6],x[5],x[4]} ,  {g[6],g[5],g[4]} , {p[6],p[5],p[4]} , G3[3] , {sum[7],sum[6],sum[5],sum[4]} ) ;
    _Psum_sparse4 _Psum_sparse4_8( {x[11],x[10],x[9],x[8]} ,  {g[10],g[9],g[8]} , {p[10],p[9],p[8]} , G3[7] , {sum[11],sum[10],sum[9],sum[8]} ) ;
    _Psum_sparse4 _Psum_sparse4_12( {x[15],x[14],x[13],x[12]} ,  {g[14],g[13],g[12]} , {p[14],p[13],p[12]} , G3[11] , {sum[15],sum[14],sum[13],sum[12]} ) ;
    _Psum_sparse4 _Psum_sparse4_16( {x[19],x[18],x[17],x[16]} ,  {g[18],g[17],g[16]} , {p[18],p[17],p[16]} , G3[15] , {sum[19],sum[18],sum[17],sum[16]} ) ;
    _Psum_sparse4 _Psum_sparse4_20( {x[23],x[22],x[21],x[20]} ,  {g[22],g[21],g[20]} , {p[22],p[21],p[20]} , G3[19] , {sum[23],sum[22],sum[21],sum[20]} ) ;
    _Psum_sparse4 _Psum_sparse4_24( {x[27],x[26],x[25],x[24]} ,  {g[26],g[25],g[24]} , {p[26],p[25],p[24]} , G3[23] , {sum[27],sum[26],sum[25],sum[24]} ) ;
    _Psum_sparse4 _Psum_sparse4_28( {x[31],x[30],x[29],x[28]} ,  {g[30],g[29],g[28]} , {p[30],p[29],p[28]} , G3[27] , {sum[31],sum[30],sum[29],sum[28]} ) ;
    _Psum_sparse4 _Psum_sparse4_32( {x[35],x[34],x[33],x[32]} ,  {g[34],g[33],g[32]} , {p[34],p[33],p[32]} , G3[31] , {sum[35],sum[34],sum[33],sum[32]} ) ;
    _Psum_sparse4 _Psum_sparse4_36( {x[39],x[38],x[37],x[36]} ,  {g[38],g[37],g[36]} , {p[38],p[37],p[36]} , G3[35] , {sum[39],sum[38],sum[37],sum[36]} ) ;
    _Psum_sparse4 _Psum_sparse4_40( {x[43],x[42],x[41],x[40]} ,  {g[42],g[41],g[40]} , {p[42],p[41],p[40]} , G3[39] , {sum[43],sum[42],sum[41],sum[40]} ) ;
    _Psum_sparse4 _Psum_sparse4_44( {x[47],x[46],x[45],x[44]} ,  {g[46],g[45],g[44]} , {p[46],p[45],p[44]} , G3[43] , {sum[47],sum[46],sum[45],sum[44]} ) ;
    _Psum_sparse4 _Psum_sparse4_48( {x[51],x[50],x[49],x[48]} ,  {g[50],g[49],g[48]} , {p[50],p[49],p[48]} , G3[47] , {sum[51],sum[50],sum[49],sum[48]} ) ;
    _Psum_sparse4 _Psum_sparse4_52( {x[55],x[54],x[53],x[52]} ,  {g[54],g[53],g[52]} , {p[54],p[53],p[52]} , G3[51] , {sum[55],sum[54],sum[53],sum[52]} ) ;
    _Psum_sparse4 _Psum_sparse4_56( {x[59],x[58],x[57],x[56]} ,  {g[58],g[57],g[56]} , {p[58],p[57],p[56]} , G3[55] , {sum[59],sum[58],sum[57],sum[56]} ) ;
    _Psum_sparse4 _Psum_sparse4_60( {x[63],x[62],x[61],x[60]} ,  {g[62],g[61],g[60]} , {p[62],p[61],p[60]} , G3[59] , {sum[63],sum[62],sum[61],sum[60]} ) ;

endmodule
