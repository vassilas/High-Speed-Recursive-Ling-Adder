// Stage 1
//--------------------------------------------------------------------------------------
module J32_stage_1(a, b, g, p, x, R1, Q1, D_r);
//
//
//
    input [31:0]a ;
    input [31:0]b ;
    output [31:0]g ;
    output [31:0]p ;
    output [31:0]x ;
    output [31:0]R1 ;
    output [31:0]Q1 ;
    output [31:0]D_r ;
    
    
    assign p[31:0] = a[31:0] | b[31:0] ;
    assign g[31:0] = a[31:0] & b[31:0] ;
    assign x[31:0] = a[31:0] ^ b[31:0] ;    
    
    assign R1[31:0] = g[31:0] | {g[30:0],g[31]};
    assign Q1[31:0] = p[31:0] & {p[30:0],p[31]} ;
    
    assign D_r[31:0] = g[31:0] | p[31:0]&{g[30:0],g[31]} | p[31:0]&{p[30:0],p[31]}&{p[29:0],p[31:30]} ;
    
endmodule


// Stage 2
//--------------------------------------------------------------------------------------
module J32_stage_2(R1, Q1, R2, Q2);
//
//
//
    input [31:0]R1;
    input [31:0]Q1;
    output [31:0]R2;
    output [31:0]Q2;

    assign R2[31:0] = R1[31:0] | {R1[29:0],R1[31:30]} | {Q1[28:0],Q1[31:29]} & {R1[27:0],R1[31:28]} | {Q1[28:0],Q1[31:29]}&{Q1[26:0],Q1[31:27]}&{R1[25:0],R1[31:26]} ;
    assign Q2[31:0] = Q1[31:0] & {Q1[29:0],Q1[31:30]} & {Q1[27:0],Q1[31:28]} & ({R1[26:0],R1[31:27]} | {Q1[25:0],Q1[31:26]});
    
endmodule



// Stage 3
//--------------------------------------------------------------------------------------
module J32_stage_3(R2, Q2, x, D_r, R3, xD);
//
//
//
    input [31:0]R2;
    input [31:0]Q2;
    input [31:0]D_r;
    input [31:0]x;
    output [31:0]R3;
    output [31:0]xD;
    
    wire [31:0]D;
    
    assign R3[31:0] = R2[31:0] | {R2[23:0],R2[31:24]} | {Q2[20:0],Q2[31:21]} & {R2[15:0],R2[31:16]} | {Q2[20:0],Q2[31:21]} & {Q2[12:0],Q2[31:13]} & {R2[7:0],R2[31:8]} ;
    
    assign D[31:0] = D_r[31:0] & ( R2[31:0] | {Q2[28:0],Q2[31:29]} ) ;
    assign xD[31:0] = x[31:0] ^ {D[30:0],D[31]} ;
    
endmodule




// Adder
//--------------------------------------------------------------------------------------
module J32_adder(a, b, sum);
//
//
//
    input [31:0]a;
    input [31:0]b;
    output [31:0]sum;
    
    wire [31:0] g ;
    wire [31:0] p ;
    wire [31:0] x ;
    wire [31:0] R1 ;
    wire [31:0] R2 ;
    wire [31:0] R3 ;
    wire [31:0] Q1 ;
    wire [31:0] Q2 ;
    wire [31:0] D_r ;
    wire [31:0] xD ;

    
    J32_stage_1 CUT1(a, b, g, p, x, R1, Q1, D_r);
    J32_stage_2 CUT2(R1, Q1, R2, Q2);
    J32_stage_3 CUT3(R2, Q2, x, D_r, R3, xD);
    

    assign sum[31:0] = ~{R3[30:0],R3[31]} & (x[31:0]) | {R3[30:0],R3[31]} & xD[31:0] ;
    
endmodule









// With D recursion Module
//------------------------------
/*
// Stage 1
//--------------------------------------------------------------------------------------
module J32D_stage_1(a, b, g, p, x, R1, Q1);
//
//
//
    input [31:0]a ;
    input [31:0]b ;
    output [31:0]g ;
    output [31:0]p ;
    output [31:0]x ;
    output [31:0]R1 ;
    output [31:0]Q1 ;

    
    
    assign p[31:0] = a[31:0] | b[31:0] ;
    assign g[31:0] = a[31:0] & b[31:0] ;
    assign x[31:0] = a[31:0] ^ b[31:0] ;    
    
    assign R1[31:0] = g[31:0] | {g[30:0],g[31]};
    assign Q1[31:0] = p[31:0] & {p[30:0],p[31]} ;
    
    
endmodule

// Stage 3
//--------------------------------------------------------------------------------------
module J32D_stage_3(R2, Q2, R3);
//
//
//
    input [31:0]R2;
    input [31:0]Q2;

    output [31:0]R3;

    

    
    assign R3[31:0] = R2[31:0] | {R2[23:0],R2[31:24]} | {Q2[20:0],Q2[31:21]} & {R2[15:0],R2[31:16]} | {Q2[20:0],Q2[31:21]} & {Q2[12:0],Q2[31:13]} & {R2[7:0],R2[31:8]} ;
    

    
endmodule


module J32_Drecursion(p, g, R2, Q2, D);
    
    input [31:0]p ;    
    input [31:0]g ;
    input [31:0]R2;
    input [31:0]Q2;

    output [31:0]D;
    
    wire [31:0]D_r;
    
    assign D_r[31:0] = g[31:0] | p[31:0]&{g[30:0],g[31]} | p[31:0]&{p[30:0],p[31]}&{p[29:0],p[31:30]} ;
    assign D[31:0] = D_r[31:0] & ( R2[31:0] | {Q2[28:0],Q2[31:29]} ) ;
     
endmodule



// Adder
//--------------------------------------------------------------------------------------
module J32_adder(a, b, sum);
//
//
//
    input [31:0]a;
    input [31:0]b;
    output [31:0]sum;
    
    wire [31:0] g ;
    wire [31:0] p ;
    wire [31:0] x ;
    wire [31:0] R1 ;
    wire [31:0] R2 ;
    wire [31:0] R3 ;
    wire [31:0] Q1 ;
    wire [31:0] Q2 ;
    wire [31:0] D ;

    
    J32D_stage_1 CUT1(a, b, g, p, x, R1, Q1);
    J32_stage_2 CUT2(R1, Q1, R2, Q2);
    J32D_stage_3 CUT3(R2, Q2, R3);
    J32_Drecursion CUT4(p, g, R2, Q2, D);

    assign sum[31:0] = ~{R3[30:0],R3[31]} & (x[31:0]) | {R3[30:0],R3[31]} & ( x[31:0] ^ {D[30:0],D[31]} ) ;
    
endmodule
*/