module P64_node_adder(a, b, sum);
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    wire [63:0]g ;
    wire [63:0]p ;
    wire [63:0]x ;
    wire [63:0]G1 ;
    wire [63:0]G2 ;
    wire [63:0]G3 ;
    wire [63:0]Pr1 ;
    wire [63:0]Pr2 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;
    _gpx _gpx_16	(a[16],	b[16],	g[16], 	p[16], 	x[16]) ;
    _gpx _gpx_17	(a[17],	b[17],	g[17], 	p[17], 	x[17]) ;
    _gpx _gpx_18	(a[18],	b[18],	g[18], 	p[18], 	x[18]) ;
    _gpx _gpx_19	(a[19],	b[19],	g[19], 	p[19], 	x[19]) ;
    _gpx _gpx_20	(a[20],	b[20],	g[20], 	p[20], 	x[20]) ;
    _gpx _gpx_21	(a[21],	b[21],	g[21], 	p[21], 	x[21]) ;
    _gpx _gpx_22	(a[22],	b[22],	g[22], 	p[22], 	x[22]) ;
    _gpx _gpx_23	(a[23],	b[23],	g[23], 	p[23], 	x[23]) ;
    _gpx _gpx_24	(a[24],	b[24],	g[24], 	p[24], 	x[24]) ;
    _gpx _gpx_25	(a[25],	b[25],	g[25], 	p[25], 	x[25]) ;
    _gpx _gpx_26	(a[26],	b[26],	g[26], 	p[26], 	x[26]) ;
    _gpx _gpx_27	(a[27],	b[27],	g[27], 	p[27], 	x[27]) ;
    _gpx _gpx_28	(a[28],	b[28],	g[28], 	p[28], 	x[28]) ;
    _gpx _gpx_29	(a[29],	b[29],	g[29], 	p[29], 	x[29]) ;
    _gpx _gpx_30	(a[30],	b[30],	g[30], 	p[30], 	x[30]) ;
    _gpx _gpx_31	(a[31],	b[31],	g[31], 	p[31], 	x[31]) ;
    _gpx _gpx_32	(a[32],	b[32],	g[32], 	p[32], 	x[32]) ;
    _gpx _gpx_33	(a[33],	b[33],	g[33], 	p[33], 	x[33]) ;
    _gpx _gpx_34	(a[34],	b[34],	g[34], 	p[34], 	x[34]) ;
    _gpx _gpx_35	(a[35],	b[35],	g[35], 	p[35], 	x[35]) ;
    _gpx _gpx_36	(a[36],	b[36],	g[36], 	p[36], 	x[36]) ;
    _gpx _gpx_37	(a[37],	b[37],	g[37], 	p[37], 	x[37]) ;
    _gpx _gpx_38	(a[38],	b[38],	g[38], 	p[38], 	x[38]) ;
    _gpx _gpx_39	(a[39],	b[39],	g[39], 	p[39], 	x[39]) ;
    _gpx _gpx_40	(a[40],	b[40],	g[40], 	p[40], 	x[40]) ;
    _gpx _gpx_41	(a[41],	b[41],	g[41], 	p[41], 	x[41]) ;
    _gpx _gpx_42	(a[42],	b[42],	g[42], 	p[42], 	x[42]) ;
    _gpx _gpx_43	(a[43],	b[43],	g[43], 	p[43], 	x[43]) ;
    _gpx _gpx_44	(a[44],	b[44],	g[44], 	p[44], 	x[44]) ;
    _gpx _gpx_45	(a[45],	b[45],	g[45], 	p[45], 	x[45]) ;
    _gpx _gpx_46	(a[46],	b[46],	g[46], 	p[46], 	x[46]) ;
    _gpx _gpx_47	(a[47],	b[47],	g[47], 	p[47], 	x[47]) ;
    _gpx _gpx_48	(a[48],	b[48],	g[48], 	p[48], 	x[48]) ;
    _gpx _gpx_49	(a[49],	b[49],	g[49], 	p[49], 	x[49]) ;
    _gpx _gpx_50	(a[50],	b[50],	g[50], 	p[50], 	x[50]) ;
    _gpx _gpx_51	(a[51],	b[51],	g[51], 	p[51], 	x[51]) ;
    _gpx _gpx_52	(a[52],	b[52],	g[52], 	p[52], 	x[52]) ;
    _gpx _gpx_53	(a[53],	b[53],	g[53], 	p[53], 	x[53]) ;
    _gpx _gpx_54	(a[54],	b[54],	g[54], 	p[54], 	x[54]) ;
    _gpx _gpx_55	(a[55],	b[55],	g[55], 	p[55], 	x[55]) ;
    _gpx _gpx_56	(a[56],	b[56],	g[56], 	p[56], 	x[56]) ;
    _gpx _gpx_57	(a[57],	b[57],	g[57], 	p[57], 	x[57]) ;
    _gpx _gpx_58	(a[58],	b[58],	g[58], 	p[58], 	x[58]) ;
    _gpx _gpx_59	(a[59],	b[59],	g[59], 	p[59], 	x[59]) ;
    _gpx _gpx_60	(a[60],	b[60],	g[60], 	p[60], 	x[60]) ;
    _gpx _gpx_61	(a[61],	b[61],	g[61], 	p[61], 	x[61]) ;
    _gpx _gpx_62	(a[62],	b[62],	g[62], 	p[62], 	x[62]) ;
    _gpx _gpx_63	(a[63],	b[63],	g[63], 	p[63], 	x[63]) ;

    _4G3P_G4 _4G3P_G4_0( {g[0],g[63],g[62],g[61]} , {p[0],p[63],p[62]} ,G1[0] ) ;
    _4G3P_G4 _4G3P_G4_1( {g[1],g[0],g[63],g[62]} , {p[1],p[0],p[63]} ,G1[1] ) ;
    _4G3P_G4 _4G3P_G4_2( {g[2],g[1],g[0],g[63]} , {p[2],p[1],p[0]} ,G1[2] ) ;
    _4G3P_G4 _4G3P_G4_3( {g[3],g[2],g[1],g[0]} , {p[3],p[2],p[1]} ,G1[3] ) ;
    _4G3P_G4 _4G3P_G4_4( {g[4],g[3],g[2],g[1]} , {p[4],p[3],p[2]} ,G1[4] ) ;
    _4G3P_G4 _4G3P_G4_5( {g[5],g[4],g[3],g[2]} , {p[5],p[4],p[3]} ,G1[5] ) ;
    _4G3P_G4 _4G3P_G4_6( {g[6],g[5],g[4],g[3]} , {p[6],p[5],p[4]} ,G1[6] ) ;
    _4G3P_G4 _4G3P_G4_7( {g[7],g[6],g[5],g[4]} , {p[7],p[6],p[5]} ,G1[7] ) ;
    _4G3P_G4 _4G3P_G4_8( {g[8],g[7],g[6],g[5]} , {p[8],p[7],p[6]} ,G1[8] ) ;
    _4G3P_G4 _4G3P_G4_9( {g[9],g[8],g[7],g[6]} , {p[9],p[8],p[7]} ,G1[9] ) ;
    _4G3P_G4 _4G3P_G4_10( {g[10],g[9],g[8],g[7]} , {p[10],p[9],p[8]} ,G1[10] ) ;
    _4G3P_G4 _4G3P_G4_11( {g[11],g[10],g[9],g[8]} , {p[11],p[10],p[9]} ,G1[11] ) ;
    _4G3P_G4 _4G3P_G4_12( {g[12],g[11],g[10],g[9]} , {p[12],p[11],p[10]} ,G1[12] ) ;
    _4G3P_G4 _4G3P_G4_13( {g[13],g[12],g[11],g[10]} , {p[13],p[12],p[11]} ,G1[13] ) ;
    _4G3P_G4 _4G3P_G4_14( {g[14],g[13],g[12],g[11]} , {p[14],p[13],p[12]} ,G1[14] ) ;
    _4G3P_G4 _4G3P_G4_15( {g[15],g[14],g[13],g[12]} , {p[15],p[14],p[13]} ,G1[15] ) ;
    _4G3P_G4 _4G3P_G4_16( {g[16],g[15],g[14],g[13]} , {p[16],p[15],p[14]} ,G1[16] ) ;
    _4G3P_G4 _4G3P_G4_17( {g[17],g[16],g[15],g[14]} , {p[17],p[16],p[15]} ,G1[17] ) ;
    _4G3P_G4 _4G3P_G4_18( {g[18],g[17],g[16],g[15]} , {p[18],p[17],p[16]} ,G1[18] ) ;
    _4G3P_G4 _4G3P_G4_19( {g[19],g[18],g[17],g[16]} , {p[19],p[18],p[17]} ,G1[19] ) ;
    _4G3P_G4 _4G3P_G4_20( {g[20],g[19],g[18],g[17]} , {p[20],p[19],p[18]} ,G1[20] ) ;
    _4G3P_G4 _4G3P_G4_21( {g[21],g[20],g[19],g[18]} , {p[21],p[20],p[19]} ,G1[21] ) ;
    _4G3P_G4 _4G3P_G4_22( {g[22],g[21],g[20],g[19]} , {p[22],p[21],p[20]} ,G1[22] ) ;
    _4G3P_G4 _4G3P_G4_23( {g[23],g[22],g[21],g[20]} , {p[23],p[22],p[21]} ,G1[23] ) ;
    _4G3P_G4 _4G3P_G4_24( {g[24],g[23],g[22],g[21]} , {p[24],p[23],p[22]} ,G1[24] ) ;
    _4G3P_G4 _4G3P_G4_25( {g[25],g[24],g[23],g[22]} , {p[25],p[24],p[23]} ,G1[25] ) ;
    _4G3P_G4 _4G3P_G4_26( {g[26],g[25],g[24],g[23]} , {p[26],p[25],p[24]} ,G1[26] ) ;
    _4G3P_G4 _4G3P_G4_27( {g[27],g[26],g[25],g[24]} , {p[27],p[26],p[25]} ,G1[27] ) ;
    _4G3P_G4 _4G3P_G4_28( {g[28],g[27],g[26],g[25]} , {p[28],p[27],p[26]} ,G1[28] ) ;
    _4G3P_G4 _4G3P_G4_29( {g[29],g[28],g[27],g[26]} , {p[29],p[28],p[27]} ,G1[29] ) ;
    _4G3P_G4 _4G3P_G4_30( {g[30],g[29],g[28],g[27]} , {p[30],p[29],p[28]} ,G1[30] ) ;
    _4G3P_G4 _4G3P_G4_31( {g[31],g[30],g[29],g[28]} , {p[31],p[30],p[29]} ,G1[31] ) ;
    _4G3P_G4 _4G3P_G4_32( {g[32],g[31],g[30],g[29]} , {p[32],p[31],p[30]} ,G1[32] ) ;
    _4G3P_G4 _4G3P_G4_33( {g[33],g[32],g[31],g[30]} , {p[33],p[32],p[31]} ,G1[33] ) ;
    _4G3P_G4 _4G3P_G4_34( {g[34],g[33],g[32],g[31]} , {p[34],p[33],p[32]} ,G1[34] ) ;
    _4G3P_G4 _4G3P_G4_35( {g[35],g[34],g[33],g[32]} , {p[35],p[34],p[33]} ,G1[35] ) ;
    _4G3P_G4 _4G3P_G4_36( {g[36],g[35],g[34],g[33]} , {p[36],p[35],p[34]} ,G1[36] ) ;
    _4G3P_G4 _4G3P_G4_37( {g[37],g[36],g[35],g[34]} , {p[37],p[36],p[35]} ,G1[37] ) ;
    _4G3P_G4 _4G3P_G4_38( {g[38],g[37],g[36],g[35]} , {p[38],p[37],p[36]} ,G1[38] ) ;
    _4G3P_G4 _4G3P_G4_39( {g[39],g[38],g[37],g[36]} , {p[39],p[38],p[37]} ,G1[39] ) ;
    _4G3P_G4 _4G3P_G4_40( {g[40],g[39],g[38],g[37]} , {p[40],p[39],p[38]} ,G1[40] ) ;
    _4G3P_G4 _4G3P_G4_41( {g[41],g[40],g[39],g[38]} , {p[41],p[40],p[39]} ,G1[41] ) ;
    _4G3P_G4 _4G3P_G4_42( {g[42],g[41],g[40],g[39]} , {p[42],p[41],p[40]} ,G1[42] ) ;
    _4G3P_G4 _4G3P_G4_43( {g[43],g[42],g[41],g[40]} , {p[43],p[42],p[41]} ,G1[43] ) ;
    _4G3P_G4 _4G3P_G4_44( {g[44],g[43],g[42],g[41]} , {p[44],p[43],p[42]} ,G1[44] ) ;
    _4G3P_G4 _4G3P_G4_45( {g[45],g[44],g[43],g[42]} , {p[45],p[44],p[43]} ,G1[45] ) ;
    _4G3P_G4 _4G3P_G4_46( {g[46],g[45],g[44],g[43]} , {p[46],p[45],p[44]} ,G1[46] ) ;
    _4G3P_G4 _4G3P_G4_47( {g[47],g[46],g[45],g[44]} , {p[47],p[46],p[45]} ,G1[47] ) ;
    _4G3P_G4 _4G3P_G4_48( {g[48],g[47],g[46],g[45]} , {p[48],p[47],p[46]} ,G1[48] ) ;
    _4G3P_G4 _4G3P_G4_49( {g[49],g[48],g[47],g[46]} , {p[49],p[48],p[47]} ,G1[49] ) ;
    _4G3P_G4 _4G3P_G4_50( {g[50],g[49],g[48],g[47]} , {p[50],p[49],p[48]} ,G1[50] ) ;
    _4G3P_G4 _4G3P_G4_51( {g[51],g[50],g[49],g[48]} , {p[51],p[50],p[49]} ,G1[51] ) ;
    _4G3P_G4 _4G3P_G4_52( {g[52],g[51],g[50],g[49]} , {p[52],p[51],p[50]} ,G1[52] ) ;
    _4G3P_G4 _4G3P_G4_53( {g[53],g[52],g[51],g[50]} , {p[53],p[52],p[51]} ,G1[53] ) ;
    _4G3P_G4 _4G3P_G4_54( {g[54],g[53],g[52],g[51]} , {p[54],p[53],p[52]} ,G1[54] ) ;
    _4G3P_G4 _4G3P_G4_55( {g[55],g[54],g[53],g[52]} , {p[55],p[54],p[53]} ,G1[55] ) ;
    _4G3P_G4 _4G3P_G4_56( {g[56],g[55],g[54],g[53]} , {p[56],p[55],p[54]} ,G1[56] ) ;
    _4G3P_G4 _4G3P_G4_57( {g[57],g[56],g[55],g[54]} , {p[57],p[56],p[55]} ,G1[57] ) ;
    _4G3P_G4 _4G3P_G4_58( {g[58],g[57],g[56],g[55]} , {p[58],p[57],p[56]} ,G1[58] ) ;
    _4G3P_G4 _4G3P_G4_59( {g[59],g[58],g[57],g[56]} , {p[59],p[58],p[57]} ,G1[59] ) ;
    _4G3P_G4 _4G3P_G4_60( {g[60],g[59],g[58],g[57]} , {p[60],p[59],p[58]} ,G1[60] ) ;
    _4G3P_G4 _4G3P_G4_61( {g[61],g[60],g[59],g[58]} , {p[61],p[60],p[59]} ,G1[61] ) ;
    _4G3P_G4 _4G3P_G4_62( {g[62],g[61],g[60],g[59]} , {p[62],p[61],p[60]} ,G1[62] ) ;
    _4G3P_G4 _4G3P_G4_63( {g[63],g[62],g[61],g[60]} , {p[63],p[62],p[61]} ,G1[63] ) ;

    _P4 _P4_0( {p[0],p[63],p[62],p[61]} ,Pr1[0] ) ;
    _P4 _P4_1( {p[1],p[0],p[63],p[62]} ,Pr1[1] ) ;
    _P4 _P4_2( {p[2],p[1],p[0],p[63]} ,Pr1[2] ) ;
    _P4 _P4_3( {p[3],p[2],p[1],p[0]} ,Pr1[3] ) ;
    _P4 _P4_4( {p[4],p[3],p[2],p[1]} ,Pr1[4] ) ;
    _P4 _P4_5( {p[5],p[4],p[3],p[2]} ,Pr1[5] ) ;
    _P4 _P4_6( {p[6],p[5],p[4],p[3]} ,Pr1[6] ) ;
    _P4 _P4_7( {p[7],p[6],p[5],p[4]} ,Pr1[7] ) ;
    _P4 _P4_8( {p[8],p[7],p[6],p[5]} ,Pr1[8] ) ;
    _P4 _P4_9( {p[9],p[8],p[7],p[6]} ,Pr1[9] ) ;
    _P4 _P4_10( {p[10],p[9],p[8],p[7]} ,Pr1[10] ) ;
    _P4 _P4_11( {p[11],p[10],p[9],p[8]} ,Pr1[11] ) ;
    _P4 _P4_12( {p[12],p[11],p[10],p[9]} ,Pr1[12] ) ;
    _P4 _P4_13( {p[13],p[12],p[11],p[10]} ,Pr1[13] ) ;
    _P4 _P4_14( {p[14],p[13],p[12],p[11]} ,Pr1[14] ) ;
    _P4 _P4_15( {p[15],p[14],p[13],p[12]} ,Pr1[15] ) ;
    _P4 _P4_16( {p[16],p[15],p[14],p[13]} ,Pr1[16] ) ;
    _P4 _P4_17( {p[17],p[16],p[15],p[14]} ,Pr1[17] ) ;
    _P4 _P4_18( {p[18],p[17],p[16],p[15]} ,Pr1[18] ) ;
    _P4 _P4_19( {p[19],p[18],p[17],p[16]} ,Pr1[19] ) ;
    _P4 _P4_20( {p[20],p[19],p[18],p[17]} ,Pr1[20] ) ;
    _P4 _P4_21( {p[21],p[20],p[19],p[18]} ,Pr1[21] ) ;
    _P4 _P4_22( {p[22],p[21],p[20],p[19]} ,Pr1[22] ) ;
    _P4 _P4_23( {p[23],p[22],p[21],p[20]} ,Pr1[23] ) ;
    _P4 _P4_24( {p[24],p[23],p[22],p[21]} ,Pr1[24] ) ;
    _P4 _P4_25( {p[25],p[24],p[23],p[22]} ,Pr1[25] ) ;
    _P4 _P4_26( {p[26],p[25],p[24],p[23]} ,Pr1[26] ) ;
    _P4 _P4_27( {p[27],p[26],p[25],p[24]} ,Pr1[27] ) ;
    _P4 _P4_28( {p[28],p[27],p[26],p[25]} ,Pr1[28] ) ;
    _P4 _P4_29( {p[29],p[28],p[27],p[26]} ,Pr1[29] ) ;
    _P4 _P4_30( {p[30],p[29],p[28],p[27]} ,Pr1[30] ) ;
    _P4 _P4_31( {p[31],p[30],p[29],p[28]} ,Pr1[31] ) ;
    _P4 _P4_32( {p[32],p[31],p[30],p[29]} ,Pr1[32] ) ;
    _P4 _P4_33( {p[33],p[32],p[31],p[30]} ,Pr1[33] ) ;
    _P4 _P4_34( {p[34],p[33],p[32],p[31]} ,Pr1[34] ) ;
    _P4 _P4_35( {p[35],p[34],p[33],p[32]} ,Pr1[35] ) ;
    _P4 _P4_36( {p[36],p[35],p[34],p[33]} ,Pr1[36] ) ;
    _P4 _P4_37( {p[37],p[36],p[35],p[34]} ,Pr1[37] ) ;
    _P4 _P4_38( {p[38],p[37],p[36],p[35]} ,Pr1[38] ) ;
    _P4 _P4_39( {p[39],p[38],p[37],p[36]} ,Pr1[39] ) ;
    _P4 _P4_40( {p[40],p[39],p[38],p[37]} ,Pr1[40] ) ;
    _P4 _P4_41( {p[41],p[40],p[39],p[38]} ,Pr1[41] ) ;
    _P4 _P4_42( {p[42],p[41],p[40],p[39]} ,Pr1[42] ) ;
    _P4 _P4_43( {p[43],p[42],p[41],p[40]} ,Pr1[43] ) ;
    _P4 _P4_44( {p[44],p[43],p[42],p[41]} ,Pr1[44] ) ;
    _P4 _P4_45( {p[45],p[44],p[43],p[42]} ,Pr1[45] ) ;
    _P4 _P4_46( {p[46],p[45],p[44],p[43]} ,Pr1[46] ) ;
    _P4 _P4_47( {p[47],p[46],p[45],p[44]} ,Pr1[47] ) ;
    _P4 _P4_48( {p[48],p[47],p[46],p[45]} ,Pr1[48] ) ;
    _P4 _P4_49( {p[49],p[48],p[47],p[46]} ,Pr1[49] ) ;
    _P4 _P4_50( {p[50],p[49],p[48],p[47]} ,Pr1[50] ) ;
    _P4 _P4_51( {p[51],p[50],p[49],p[48]} ,Pr1[51] ) ;
    _P4 _P4_52( {p[52],p[51],p[50],p[49]} ,Pr1[52] ) ;
    _P4 _P4_53( {p[53],p[52],p[51],p[50]} ,Pr1[53] ) ;
    _P4 _P4_54( {p[54],p[53],p[52],p[51]} ,Pr1[54] ) ;
    _P4 _P4_55( {p[55],p[54],p[53],p[52]} ,Pr1[55] ) ;
    _P4 _P4_56( {p[56],p[55],p[54],p[53]} ,Pr1[56] ) ;
    _P4 _P4_57( {p[57],p[56],p[55],p[54]} ,Pr1[57] ) ;
    _P4 _P4_58( {p[58],p[57],p[56],p[55]} ,Pr1[58] ) ;
    _P4 _P4_59( {p[59],p[58],p[57],p[56]} ,Pr1[59] ) ;
    _P4 _P4_60( {p[60],p[59],p[58],p[57]} ,Pr1[60] ) ;
    _P4 _P4_61( {p[61],p[60],p[59],p[58]} ,Pr1[61] ) ;
    _P4 _P4_62( {p[62],p[61],p[60],p[59]} ,Pr1[62] ) ;
    _P4 _P4_63( {p[63],p[62],p[61],p[60]} ,Pr1[63] ) ;

    _4G3P_G4 _4G3P_G4_64( {G1[0],G1[60],G1[56],G1[52]} , {Pr1[0],Pr1[60],Pr1[56]} ,G2[0] ) ;
    _4G3P_G4 _4G3P_G4_65( {G1[1],G1[61],G1[57],G1[53]} , {Pr1[1],Pr1[61],Pr1[57]} ,G2[1] ) ;
    _4G3P_G4 _4G3P_G4_66( {G1[2],G1[62],G1[58],G1[54]} , {Pr1[2],Pr1[62],Pr1[58]} ,G2[2] ) ;
    _4G3P_G4 _4G3P_G4_67( {G1[3],G1[63],G1[59],G1[55]} , {Pr1[3],Pr1[63],Pr1[59]} ,G2[3] ) ;
    _4G3P_G4 _4G3P_G4_68( {G1[4],G1[0],G1[60],G1[56]} , {Pr1[4],Pr1[0],Pr1[60]} ,G2[4] ) ;
    _4G3P_G4 _4G3P_G4_69( {G1[5],G1[1],G1[61],G1[57]} , {Pr1[5],Pr1[1],Pr1[61]} ,G2[5] ) ;
    _4G3P_G4 _4G3P_G4_70( {G1[6],G1[2],G1[62],G1[58]} , {Pr1[6],Pr1[2],Pr1[62]} ,G2[6] ) ;
    _4G3P_G4 _4G3P_G4_71( {G1[7],G1[3],G1[63],G1[59]} , {Pr1[7],Pr1[3],Pr1[63]} ,G2[7] ) ;
    _4G3P_G4 _4G3P_G4_72( {G1[8],G1[4],G1[0],G1[60]} , {Pr1[8],Pr1[4],Pr1[0]} ,G2[8] ) ;
    _4G3P_G4 _4G3P_G4_73( {G1[9],G1[5],G1[1],G1[61]} , {Pr1[9],Pr1[5],Pr1[1]} ,G2[9] ) ;
    _4G3P_G4 _4G3P_G4_74( {G1[10],G1[6],G1[2],G1[62]} , {Pr1[10],Pr1[6],Pr1[2]} ,G2[10] ) ;
    _4G3P_G4 _4G3P_G4_75( {G1[11],G1[7],G1[3],G1[63]} , {Pr1[11],Pr1[7],Pr1[3]} ,G2[11] ) ;
    _4G3P_G4 _4G3P_G4_76( {G1[12],G1[8],G1[4],G1[0]} , {Pr1[12],Pr1[8],Pr1[4]} ,G2[12] ) ;
    _4G3P_G4 _4G3P_G4_77( {G1[13],G1[9],G1[5],G1[1]} , {Pr1[13],Pr1[9],Pr1[5]} ,G2[13] ) ;
    _4G3P_G4 _4G3P_G4_78( {G1[14],G1[10],G1[6],G1[2]} , {Pr1[14],Pr1[10],Pr1[6]} ,G2[14] ) ;
    _4G3P_G4 _4G3P_G4_79( {G1[15],G1[11],G1[7],G1[3]} , {Pr1[15],Pr1[11],Pr1[7]} ,G2[15] ) ;
    _4G3P_G4 _4G3P_G4_80( {G1[16],G1[12],G1[8],G1[4]} , {Pr1[16],Pr1[12],Pr1[8]} ,G2[16] ) ;
    _4G3P_G4 _4G3P_G4_81( {G1[17],G1[13],G1[9],G1[5]} , {Pr1[17],Pr1[13],Pr1[9]} ,G2[17] ) ;
    _4G3P_G4 _4G3P_G4_82( {G1[18],G1[14],G1[10],G1[6]} , {Pr1[18],Pr1[14],Pr1[10]} ,G2[18] ) ;
    _4G3P_G4 _4G3P_G4_83( {G1[19],G1[15],G1[11],G1[7]} , {Pr1[19],Pr1[15],Pr1[11]} ,G2[19] ) ;
    _4G3P_G4 _4G3P_G4_84( {G1[20],G1[16],G1[12],G1[8]} , {Pr1[20],Pr1[16],Pr1[12]} ,G2[20] ) ;
    _4G3P_G4 _4G3P_G4_85( {G1[21],G1[17],G1[13],G1[9]} , {Pr1[21],Pr1[17],Pr1[13]} ,G2[21] ) ;
    _4G3P_G4 _4G3P_G4_86( {G1[22],G1[18],G1[14],G1[10]} , {Pr1[22],Pr1[18],Pr1[14]} ,G2[22] ) ;
    _4G3P_G4 _4G3P_G4_87( {G1[23],G1[19],G1[15],G1[11]} , {Pr1[23],Pr1[19],Pr1[15]} ,G2[23] ) ;
    _4G3P_G4 _4G3P_G4_88( {G1[24],G1[20],G1[16],G1[12]} , {Pr1[24],Pr1[20],Pr1[16]} ,G2[24] ) ;
    _4G3P_G4 _4G3P_G4_89( {G1[25],G1[21],G1[17],G1[13]} , {Pr1[25],Pr1[21],Pr1[17]} ,G2[25] ) ;
    _4G3P_G4 _4G3P_G4_90( {G1[26],G1[22],G1[18],G1[14]} , {Pr1[26],Pr1[22],Pr1[18]} ,G2[26] ) ;
    _4G3P_G4 _4G3P_G4_91( {G1[27],G1[23],G1[19],G1[15]} , {Pr1[27],Pr1[23],Pr1[19]} ,G2[27] ) ;
    _4G3P_G4 _4G3P_G4_92( {G1[28],G1[24],G1[20],G1[16]} , {Pr1[28],Pr1[24],Pr1[20]} ,G2[28] ) ;
    _4G3P_G4 _4G3P_G4_93( {G1[29],G1[25],G1[21],G1[17]} , {Pr1[29],Pr1[25],Pr1[21]} ,G2[29] ) ;
    _4G3P_G4 _4G3P_G4_94( {G1[30],G1[26],G1[22],G1[18]} , {Pr1[30],Pr1[26],Pr1[22]} ,G2[30] ) ;
    _4G3P_G4 _4G3P_G4_95( {G1[31],G1[27],G1[23],G1[19]} , {Pr1[31],Pr1[27],Pr1[23]} ,G2[31] ) ;
    _4G3P_G4 _4G3P_G4_96( {G1[32],G1[28],G1[24],G1[20]} , {Pr1[32],Pr1[28],Pr1[24]} ,G2[32] ) ;
    _4G3P_G4 _4G3P_G4_97( {G1[33],G1[29],G1[25],G1[21]} , {Pr1[33],Pr1[29],Pr1[25]} ,G2[33] ) ;
    _4G3P_G4 _4G3P_G4_98( {G1[34],G1[30],G1[26],G1[22]} , {Pr1[34],Pr1[30],Pr1[26]} ,G2[34] ) ;
    _4G3P_G4 _4G3P_G4_99( {G1[35],G1[31],G1[27],G1[23]} , {Pr1[35],Pr1[31],Pr1[27]} ,G2[35] ) ;
    _4G3P_G4 _4G3P_G4_100( {G1[36],G1[32],G1[28],G1[24]} , {Pr1[36],Pr1[32],Pr1[28]} ,G2[36] ) ;
    _4G3P_G4 _4G3P_G4_101( {G1[37],G1[33],G1[29],G1[25]} , {Pr1[37],Pr1[33],Pr1[29]} ,G2[37] ) ;
    _4G3P_G4 _4G3P_G4_102( {G1[38],G1[34],G1[30],G1[26]} , {Pr1[38],Pr1[34],Pr1[30]} ,G2[38] ) ;
    _4G3P_G4 _4G3P_G4_103( {G1[39],G1[35],G1[31],G1[27]} , {Pr1[39],Pr1[35],Pr1[31]} ,G2[39] ) ;
    _4G3P_G4 _4G3P_G4_104( {G1[40],G1[36],G1[32],G1[28]} , {Pr1[40],Pr1[36],Pr1[32]} ,G2[40] ) ;
    _4G3P_G4 _4G3P_G4_105( {G1[41],G1[37],G1[33],G1[29]} , {Pr1[41],Pr1[37],Pr1[33]} ,G2[41] ) ;
    _4G3P_G4 _4G3P_G4_106( {G1[42],G1[38],G1[34],G1[30]} , {Pr1[42],Pr1[38],Pr1[34]} ,G2[42] ) ;
    _4G3P_G4 _4G3P_G4_107( {G1[43],G1[39],G1[35],G1[31]} , {Pr1[43],Pr1[39],Pr1[35]} ,G2[43] ) ;
    _4G3P_G4 _4G3P_G4_108( {G1[44],G1[40],G1[36],G1[32]} , {Pr1[44],Pr1[40],Pr1[36]} ,G2[44] ) ;
    _4G3P_G4 _4G3P_G4_109( {G1[45],G1[41],G1[37],G1[33]} , {Pr1[45],Pr1[41],Pr1[37]} ,G2[45] ) ;
    _4G3P_G4 _4G3P_G4_110( {G1[46],G1[42],G1[38],G1[34]} , {Pr1[46],Pr1[42],Pr1[38]} ,G2[46] ) ;
    _4G3P_G4 _4G3P_G4_111( {G1[47],G1[43],G1[39],G1[35]} , {Pr1[47],Pr1[43],Pr1[39]} ,G2[47] ) ;
    _4G3P_G4 _4G3P_G4_112( {G1[48],G1[44],G1[40],G1[36]} , {Pr1[48],Pr1[44],Pr1[40]} ,G2[48] ) ;
    _4G3P_G4 _4G3P_G4_113( {G1[49],G1[45],G1[41],G1[37]} , {Pr1[49],Pr1[45],Pr1[41]} ,G2[49] ) ;
    _4G3P_G4 _4G3P_G4_114( {G1[50],G1[46],G1[42],G1[38]} , {Pr1[50],Pr1[46],Pr1[42]} ,G2[50] ) ;
    _4G3P_G4 _4G3P_G4_115( {G1[51],G1[47],G1[43],G1[39]} , {Pr1[51],Pr1[47],Pr1[43]} ,G2[51] ) ;
    _4G3P_G4 _4G3P_G4_116( {G1[52],G1[48],G1[44],G1[40]} , {Pr1[52],Pr1[48],Pr1[44]} ,G2[52] ) ;
    _4G3P_G4 _4G3P_G4_117( {G1[53],G1[49],G1[45],G1[41]} , {Pr1[53],Pr1[49],Pr1[45]} ,G2[53] ) ;
    _4G3P_G4 _4G3P_G4_118( {G1[54],G1[50],G1[46],G1[42]} , {Pr1[54],Pr1[50],Pr1[46]} ,G2[54] ) ;
    _4G3P_G4 _4G3P_G4_119( {G1[55],G1[51],G1[47],G1[43]} , {Pr1[55],Pr1[51],Pr1[47]} ,G2[55] ) ;
    _4G3P_G4 _4G3P_G4_120( {G1[56],G1[52],G1[48],G1[44]} , {Pr1[56],Pr1[52],Pr1[48]} ,G2[56] ) ;
    _4G3P_G4 _4G3P_G4_121( {G1[57],G1[53],G1[49],G1[45]} , {Pr1[57],Pr1[53],Pr1[49]} ,G2[57] ) ;
    _4G3P_G4 _4G3P_G4_122( {G1[58],G1[54],G1[50],G1[46]} , {Pr1[58],Pr1[54],Pr1[50]} ,G2[58] ) ;
    _4G3P_G4 _4G3P_G4_123( {G1[59],G1[55],G1[51],G1[47]} , {Pr1[59],Pr1[55],Pr1[51]} ,G2[59] ) ;
    _4G3P_G4 _4G3P_G4_124( {G1[60],G1[56],G1[52],G1[48]} , {Pr1[60],Pr1[56],Pr1[52]} ,G2[60] ) ;
    _4G3P_G4 _4G3P_G4_125( {G1[61],G1[57],G1[53],G1[49]} , {Pr1[61],Pr1[57],Pr1[53]} ,G2[61] ) ;
    _4G3P_G4 _4G3P_G4_126( {G1[62],G1[58],G1[54],G1[50]} , {Pr1[62],Pr1[58],Pr1[54]} ,G2[62] ) ;
    _4G3P_G4 _4G3P_G4_127( {G1[63],G1[59],G1[55],G1[51]} , {Pr1[63],Pr1[59],Pr1[55]} ,G2[63] ) ;

    _P4 _P4_64( {Pr1[0],Pr1[60],Pr1[56],Pr1[52]} ,Pr2[0] ) ;
    _P4 _P4_65( {Pr1[1],Pr1[61],Pr1[57],Pr1[53]} ,Pr2[1] ) ;
    _P4 _P4_66( {Pr1[2],Pr1[62],Pr1[58],Pr1[54]} ,Pr2[2] ) ;
    _P4 _P4_67( {Pr1[3],Pr1[63],Pr1[59],Pr1[55]} ,Pr2[3] ) ;
    _P4 _P4_68( {Pr1[4],Pr1[0],Pr1[60],Pr1[56]} ,Pr2[4] ) ;
    _P4 _P4_69( {Pr1[5],Pr1[1],Pr1[61],Pr1[57]} ,Pr2[5] ) ;
    _P4 _P4_70( {Pr1[6],Pr1[2],Pr1[62],Pr1[58]} ,Pr2[6] ) ;
    _P4 _P4_71( {Pr1[7],Pr1[3],Pr1[63],Pr1[59]} ,Pr2[7] ) ;
    _P4 _P4_72( {Pr1[8],Pr1[4],Pr1[0],Pr1[60]} ,Pr2[8] ) ;
    _P4 _P4_73( {Pr1[9],Pr1[5],Pr1[1],Pr1[61]} ,Pr2[9] ) ;
    _P4 _P4_74( {Pr1[10],Pr1[6],Pr1[2],Pr1[62]} ,Pr2[10] ) ;
    _P4 _P4_75( {Pr1[11],Pr1[7],Pr1[3],Pr1[63]} ,Pr2[11] ) ;
    _P4 _P4_76( {Pr1[12],Pr1[8],Pr1[4],Pr1[0]} ,Pr2[12] ) ;
    _P4 _P4_77( {Pr1[13],Pr1[9],Pr1[5],Pr1[1]} ,Pr2[13] ) ;
    _P4 _P4_78( {Pr1[14],Pr1[10],Pr1[6],Pr1[2]} ,Pr2[14] ) ;
    _P4 _P4_79( {Pr1[15],Pr1[11],Pr1[7],Pr1[3]} ,Pr2[15] ) ;
    _P4 _P4_80( {Pr1[16],Pr1[12],Pr1[8],Pr1[4]} ,Pr2[16] ) ;
    _P4 _P4_81( {Pr1[17],Pr1[13],Pr1[9],Pr1[5]} ,Pr2[17] ) ;
    _P4 _P4_82( {Pr1[18],Pr1[14],Pr1[10],Pr1[6]} ,Pr2[18] ) ;
    _P4 _P4_83( {Pr1[19],Pr1[15],Pr1[11],Pr1[7]} ,Pr2[19] ) ;
    _P4 _P4_84( {Pr1[20],Pr1[16],Pr1[12],Pr1[8]} ,Pr2[20] ) ;
    _P4 _P4_85( {Pr1[21],Pr1[17],Pr1[13],Pr1[9]} ,Pr2[21] ) ;
    _P4 _P4_86( {Pr1[22],Pr1[18],Pr1[14],Pr1[10]} ,Pr2[22] ) ;
    _P4 _P4_87( {Pr1[23],Pr1[19],Pr1[15],Pr1[11]} ,Pr2[23] ) ;
    _P4 _P4_88( {Pr1[24],Pr1[20],Pr1[16],Pr1[12]} ,Pr2[24] ) ;
    _P4 _P4_89( {Pr1[25],Pr1[21],Pr1[17],Pr1[13]} ,Pr2[25] ) ;
    _P4 _P4_90( {Pr1[26],Pr1[22],Pr1[18],Pr1[14]} ,Pr2[26] ) ;
    _P4 _P4_91( {Pr1[27],Pr1[23],Pr1[19],Pr1[15]} ,Pr2[27] ) ;
    _P4 _P4_92( {Pr1[28],Pr1[24],Pr1[20],Pr1[16]} ,Pr2[28] ) ;
    _P4 _P4_93( {Pr1[29],Pr1[25],Pr1[21],Pr1[17]} ,Pr2[29] ) ;
    _P4 _P4_94( {Pr1[30],Pr1[26],Pr1[22],Pr1[18]} ,Pr2[30] ) ;
    _P4 _P4_95( {Pr1[31],Pr1[27],Pr1[23],Pr1[19]} ,Pr2[31] ) ;
    _P4 _P4_96( {Pr1[32],Pr1[28],Pr1[24],Pr1[20]} ,Pr2[32] ) ;
    _P4 _P4_97( {Pr1[33],Pr1[29],Pr1[25],Pr1[21]} ,Pr2[33] ) ;
    _P4 _P4_98( {Pr1[34],Pr1[30],Pr1[26],Pr1[22]} ,Pr2[34] ) ;
    _P4 _P4_99( {Pr1[35],Pr1[31],Pr1[27],Pr1[23]} ,Pr2[35] ) ;
    _P4 _P4_100( {Pr1[36],Pr1[32],Pr1[28],Pr1[24]} ,Pr2[36] ) ;
    _P4 _P4_101( {Pr1[37],Pr1[33],Pr1[29],Pr1[25]} ,Pr2[37] ) ;
    _P4 _P4_102( {Pr1[38],Pr1[34],Pr1[30],Pr1[26]} ,Pr2[38] ) ;
    _P4 _P4_103( {Pr1[39],Pr1[35],Pr1[31],Pr1[27]} ,Pr2[39] ) ;
    _P4 _P4_104( {Pr1[40],Pr1[36],Pr1[32],Pr1[28]} ,Pr2[40] ) ;
    _P4 _P4_105( {Pr1[41],Pr1[37],Pr1[33],Pr1[29]} ,Pr2[41] ) ;
    _P4 _P4_106( {Pr1[42],Pr1[38],Pr1[34],Pr1[30]} ,Pr2[42] ) ;
    _P4 _P4_107( {Pr1[43],Pr1[39],Pr1[35],Pr1[31]} ,Pr2[43] ) ;
    _P4 _P4_108( {Pr1[44],Pr1[40],Pr1[36],Pr1[32]} ,Pr2[44] ) ;
    _P4 _P4_109( {Pr1[45],Pr1[41],Pr1[37],Pr1[33]} ,Pr2[45] ) ;
    _P4 _P4_110( {Pr1[46],Pr1[42],Pr1[38],Pr1[34]} ,Pr2[46] ) ;
    _P4 _P4_111( {Pr1[47],Pr1[43],Pr1[39],Pr1[35]} ,Pr2[47] ) ;
    _P4 _P4_112( {Pr1[48],Pr1[44],Pr1[40],Pr1[36]} ,Pr2[48] ) ;
    _P4 _P4_113( {Pr1[49],Pr1[45],Pr1[41],Pr1[37]} ,Pr2[49] ) ;
    _P4 _P4_114( {Pr1[50],Pr1[46],Pr1[42],Pr1[38]} ,Pr2[50] ) ;
    _P4 _P4_115( {Pr1[51],Pr1[47],Pr1[43],Pr1[39]} ,Pr2[51] ) ;
    _P4 _P4_116( {Pr1[52],Pr1[48],Pr1[44],Pr1[40]} ,Pr2[52] ) ;
    _P4 _P4_117( {Pr1[53],Pr1[49],Pr1[45],Pr1[41]} ,Pr2[53] ) ;
    _P4 _P4_118( {Pr1[54],Pr1[50],Pr1[46],Pr1[42]} ,Pr2[54] ) ;
    _P4 _P4_119( {Pr1[55],Pr1[51],Pr1[47],Pr1[43]} ,Pr2[55] ) ;
    _P4 _P4_120( {Pr1[56],Pr1[52],Pr1[48],Pr1[44]} ,Pr2[56] ) ;
    _P4 _P4_121( {Pr1[57],Pr1[53],Pr1[49],Pr1[45]} ,Pr2[57] ) ;
    _P4 _P4_122( {Pr1[58],Pr1[54],Pr1[50],Pr1[46]} ,Pr2[58] ) ;
    _P4 _P4_123( {Pr1[59],Pr1[55],Pr1[51],Pr1[47]} ,Pr2[59] ) ;
    _P4 _P4_124( {Pr1[60],Pr1[56],Pr1[52],Pr1[48]} ,Pr2[60] ) ;
    _P4 _P4_125( {Pr1[61],Pr1[57],Pr1[53],Pr1[49]} ,Pr2[61] ) ;
    _P4 _P4_126( {Pr1[62],Pr1[58],Pr1[54],Pr1[50]} ,Pr2[62] ) ;
    _P4 _P4_127( {Pr1[63],Pr1[59],Pr1[55],Pr1[51]} ,Pr2[63] ) ;

    _4G3P_G4 _4G3P_G4_128( {G2[0],G2[48],G2[32],G2[16]} , {Pr2[0],Pr2[48],Pr2[32]} ,G3[0] ) ;
    _4G3P_G4 _4G3P_G4_129( {G2[1],G2[49],G2[33],G2[17]} , {Pr2[1],Pr2[49],Pr2[33]} ,G3[1] ) ;
    _4G3P_G4 _4G3P_G4_130( {G2[2],G2[50],G2[34],G2[18]} , {Pr2[2],Pr2[50],Pr2[34]} ,G3[2] ) ;
    _4G3P_G4 _4G3P_G4_131( {G2[3],G2[51],G2[35],G2[19]} , {Pr2[3],Pr2[51],Pr2[35]} ,G3[3] ) ;
    _4G3P_G4 _4G3P_G4_132( {G2[4],G2[52],G2[36],G2[20]} , {Pr2[4],Pr2[52],Pr2[36]} ,G3[4] ) ;
    _4G3P_G4 _4G3P_G4_133( {G2[5],G2[53],G2[37],G2[21]} , {Pr2[5],Pr2[53],Pr2[37]} ,G3[5] ) ;
    _4G3P_G4 _4G3P_G4_134( {G2[6],G2[54],G2[38],G2[22]} , {Pr2[6],Pr2[54],Pr2[38]} ,G3[6] ) ;
    _4G3P_G4 _4G3P_G4_135( {G2[7],G2[55],G2[39],G2[23]} , {Pr2[7],Pr2[55],Pr2[39]} ,G3[7] ) ;
    _4G3P_G4 _4G3P_G4_136( {G2[8],G2[56],G2[40],G2[24]} , {Pr2[8],Pr2[56],Pr2[40]} ,G3[8] ) ;
    _4G3P_G4 _4G3P_G4_137( {G2[9],G2[57],G2[41],G2[25]} , {Pr2[9],Pr2[57],Pr2[41]} ,G3[9] ) ;
    _4G3P_G4 _4G3P_G4_138( {G2[10],G2[58],G2[42],G2[26]} , {Pr2[10],Pr2[58],Pr2[42]} ,G3[10] ) ;
    _4G3P_G4 _4G3P_G4_139( {G2[11],G2[59],G2[43],G2[27]} , {Pr2[11],Pr2[59],Pr2[43]} ,G3[11] ) ;
    _4G3P_G4 _4G3P_G4_140( {G2[12],G2[60],G2[44],G2[28]} , {Pr2[12],Pr2[60],Pr2[44]} ,G3[12] ) ;
    _4G3P_G4 _4G3P_G4_141( {G2[13],G2[61],G2[45],G2[29]} , {Pr2[13],Pr2[61],Pr2[45]} ,G3[13] ) ;
    _4G3P_G4 _4G3P_G4_142( {G2[14],G2[62],G2[46],G2[30]} , {Pr2[14],Pr2[62],Pr2[46]} ,G3[14] ) ;
    _4G3P_G4 _4G3P_G4_143( {G2[15],G2[63],G2[47],G2[31]} , {Pr2[15],Pr2[63],Pr2[47]} ,G3[15] ) ;
    _4G3P_G4 _4G3P_G4_144( {G2[16],G2[0],G2[48],G2[32]} , {Pr2[16],Pr2[0],Pr2[48]} ,G3[16] ) ;
    _4G3P_G4 _4G3P_G4_145( {G2[17],G2[1],G2[49],G2[33]} , {Pr2[17],Pr2[1],Pr2[49]} ,G3[17] ) ;
    _4G3P_G4 _4G3P_G4_146( {G2[18],G2[2],G2[50],G2[34]} , {Pr2[18],Pr2[2],Pr2[50]} ,G3[18] ) ;
    _4G3P_G4 _4G3P_G4_147( {G2[19],G2[3],G2[51],G2[35]} , {Pr2[19],Pr2[3],Pr2[51]} ,G3[19] ) ;
    _4G3P_G4 _4G3P_G4_148( {G2[20],G2[4],G2[52],G2[36]} , {Pr2[20],Pr2[4],Pr2[52]} ,G3[20] ) ;
    _4G3P_G4 _4G3P_G4_149( {G2[21],G2[5],G2[53],G2[37]} , {Pr2[21],Pr2[5],Pr2[53]} ,G3[21] ) ;
    _4G3P_G4 _4G3P_G4_150( {G2[22],G2[6],G2[54],G2[38]} , {Pr2[22],Pr2[6],Pr2[54]} ,G3[22] ) ;
    _4G3P_G4 _4G3P_G4_151( {G2[23],G2[7],G2[55],G2[39]} , {Pr2[23],Pr2[7],Pr2[55]} ,G3[23] ) ;
    _4G3P_G4 _4G3P_G4_152( {G2[24],G2[8],G2[56],G2[40]} , {Pr2[24],Pr2[8],Pr2[56]} ,G3[24] ) ;
    _4G3P_G4 _4G3P_G4_153( {G2[25],G2[9],G2[57],G2[41]} , {Pr2[25],Pr2[9],Pr2[57]} ,G3[25] ) ;
    _4G3P_G4 _4G3P_G4_154( {G2[26],G2[10],G2[58],G2[42]} , {Pr2[26],Pr2[10],Pr2[58]} ,G3[26] ) ;
    _4G3P_G4 _4G3P_G4_155( {G2[27],G2[11],G2[59],G2[43]} , {Pr2[27],Pr2[11],Pr2[59]} ,G3[27] ) ;
    _4G3P_G4 _4G3P_G4_156( {G2[28],G2[12],G2[60],G2[44]} , {Pr2[28],Pr2[12],Pr2[60]} ,G3[28] ) ;
    _4G3P_G4 _4G3P_G4_157( {G2[29],G2[13],G2[61],G2[45]} , {Pr2[29],Pr2[13],Pr2[61]} ,G3[29] ) ;
    _4G3P_G4 _4G3P_G4_158( {G2[30],G2[14],G2[62],G2[46]} , {Pr2[30],Pr2[14],Pr2[62]} ,G3[30] ) ;
    _4G3P_G4 _4G3P_G4_159( {G2[31],G2[15],G2[63],G2[47]} , {Pr2[31],Pr2[15],Pr2[63]} ,G3[31] ) ;
    _4G3P_G4 _4G3P_G4_160( {G2[32],G2[16],G2[0],G2[48]} , {Pr2[32],Pr2[16],Pr2[0]} ,G3[32] ) ;
    _4G3P_G4 _4G3P_G4_161( {G2[33],G2[17],G2[1],G2[49]} , {Pr2[33],Pr2[17],Pr2[1]} ,G3[33] ) ;
    _4G3P_G4 _4G3P_G4_162( {G2[34],G2[18],G2[2],G2[50]} , {Pr2[34],Pr2[18],Pr2[2]} ,G3[34] ) ;
    _4G3P_G4 _4G3P_G4_163( {G2[35],G2[19],G2[3],G2[51]} , {Pr2[35],Pr2[19],Pr2[3]} ,G3[35] ) ;
    _4G3P_G4 _4G3P_G4_164( {G2[36],G2[20],G2[4],G2[52]} , {Pr2[36],Pr2[20],Pr2[4]} ,G3[36] ) ;
    _4G3P_G4 _4G3P_G4_165( {G2[37],G2[21],G2[5],G2[53]} , {Pr2[37],Pr2[21],Pr2[5]} ,G3[37] ) ;
    _4G3P_G4 _4G3P_G4_166( {G2[38],G2[22],G2[6],G2[54]} , {Pr2[38],Pr2[22],Pr2[6]} ,G3[38] ) ;
    _4G3P_G4 _4G3P_G4_167( {G2[39],G2[23],G2[7],G2[55]} , {Pr2[39],Pr2[23],Pr2[7]} ,G3[39] ) ;
    _4G3P_G4 _4G3P_G4_168( {G2[40],G2[24],G2[8],G2[56]} , {Pr2[40],Pr2[24],Pr2[8]} ,G3[40] ) ;
    _4G3P_G4 _4G3P_G4_169( {G2[41],G2[25],G2[9],G2[57]} , {Pr2[41],Pr2[25],Pr2[9]} ,G3[41] ) ;
    _4G3P_G4 _4G3P_G4_170( {G2[42],G2[26],G2[10],G2[58]} , {Pr2[42],Pr2[26],Pr2[10]} ,G3[42] ) ;
    _4G3P_G4 _4G3P_G4_171( {G2[43],G2[27],G2[11],G2[59]} , {Pr2[43],Pr2[27],Pr2[11]} ,G3[43] ) ;
    _4G3P_G4 _4G3P_G4_172( {G2[44],G2[28],G2[12],G2[60]} , {Pr2[44],Pr2[28],Pr2[12]} ,G3[44] ) ;
    _4G3P_G4 _4G3P_G4_173( {G2[45],G2[29],G2[13],G2[61]} , {Pr2[45],Pr2[29],Pr2[13]} ,G3[45] ) ;
    _4G3P_G4 _4G3P_G4_174( {G2[46],G2[30],G2[14],G2[62]} , {Pr2[46],Pr2[30],Pr2[14]} ,G3[46] ) ;
    _4G3P_G4 _4G3P_G4_175( {G2[47],G2[31],G2[15],G2[63]} , {Pr2[47],Pr2[31],Pr2[15]} ,G3[47] ) ;
    _4G3P_G4 _4G3P_G4_176( {G2[48],G2[32],G2[16],G2[0]} , {Pr2[48],Pr2[32],Pr2[16]} ,G3[48] ) ;
    _4G3P_G4 _4G3P_G4_177( {G2[49],G2[33],G2[17],G2[1]} , {Pr2[49],Pr2[33],Pr2[17]} ,G3[49] ) ;
    _4G3P_G4 _4G3P_G4_178( {G2[50],G2[34],G2[18],G2[2]} , {Pr2[50],Pr2[34],Pr2[18]} ,G3[50] ) ;
    _4G3P_G4 _4G3P_G4_179( {G2[51],G2[35],G2[19],G2[3]} , {Pr2[51],Pr2[35],Pr2[19]} ,G3[51] ) ;
    _4G3P_G4 _4G3P_G4_180( {G2[52],G2[36],G2[20],G2[4]} , {Pr2[52],Pr2[36],Pr2[20]} ,G3[52] ) ;
    _4G3P_G4 _4G3P_G4_181( {G2[53],G2[37],G2[21],G2[5]} , {Pr2[53],Pr2[37],Pr2[21]} ,G3[53] ) ;
    _4G3P_G4 _4G3P_G4_182( {G2[54],G2[38],G2[22],G2[6]} , {Pr2[54],Pr2[38],Pr2[22]} ,G3[54] ) ;
    _4G3P_G4 _4G3P_G4_183( {G2[55],G2[39],G2[23],G2[7]} , {Pr2[55],Pr2[39],Pr2[23]} ,G3[55] ) ;
    _4G3P_G4 _4G3P_G4_184( {G2[56],G2[40],G2[24],G2[8]} , {Pr2[56],Pr2[40],Pr2[24]} ,G3[56] ) ;
    _4G3P_G4 _4G3P_G4_185( {G2[57],G2[41],G2[25],G2[9]} , {Pr2[57],Pr2[41],Pr2[25]} ,G3[57] ) ;
    _4G3P_G4 _4G3P_G4_186( {G2[58],G2[42],G2[26],G2[10]} , {Pr2[58],Pr2[42],Pr2[26]} ,G3[58] ) ;
    _4G3P_G4 _4G3P_G4_187( {G2[59],G2[43],G2[27],G2[11]} , {Pr2[59],Pr2[43],Pr2[27]} ,G3[59] ) ;
    _4G3P_G4 _4G3P_G4_188( {G2[60],G2[44],G2[28],G2[12]} , {Pr2[60],Pr2[44],Pr2[28]} ,G3[60] ) ;
    _4G3P_G4 _4G3P_G4_189( {G2[61],G2[45],G2[29],G2[13]} , {Pr2[61],Pr2[45],Pr2[29]} ,G3[61] ) ;
    _4G3P_G4 _4G3P_G4_190( {G2[62],G2[46],G2[30],G2[14]} , {Pr2[62],Pr2[46],Pr2[30]} ,G3[62] ) ;
    _4G3P_G4 _4G3P_G4_191( {G2[63],G2[47],G2[31],G2[15]} , {Pr2[63],Pr2[47],Pr2[31]} ,G3[63] ) ;

    _Psum _Psum_0( x[0] , G3[63] , sum[0] ) ;
    _Psum _Psum_1( x[1] , G3[0] , sum[1] ) ;
    _Psum _Psum_2( x[2] , G3[1] , sum[2] ) ;
    _Psum _Psum_3( x[3] , G3[2] , sum[3] ) ;
    _Psum _Psum_4( x[4] , G3[3] , sum[4] ) ;
    _Psum _Psum_5( x[5] , G3[4] , sum[5] ) ;
    _Psum _Psum_6( x[6] , G3[5] , sum[6] ) ;
    _Psum _Psum_7( x[7] , G3[6] , sum[7] ) ;
    _Psum _Psum_8( x[8] , G3[7] , sum[8] ) ;
    _Psum _Psum_9( x[9] , G3[8] , sum[9] ) ;
    _Psum _Psum_10( x[10] , G3[9] , sum[10] ) ;
    _Psum _Psum_11( x[11] , G3[10] , sum[11] ) ;
    _Psum _Psum_12( x[12] , G3[11] , sum[12] ) ;
    _Psum _Psum_13( x[13] , G3[12] , sum[13] ) ;
    _Psum _Psum_14( x[14] , G3[13] , sum[14] ) ;
    _Psum _Psum_15( x[15] , G3[14] , sum[15] ) ;
    _Psum _Psum_16( x[16] , G3[15] , sum[16] ) ;
    _Psum _Psum_17( x[17] , G3[16] , sum[17] ) ;
    _Psum _Psum_18( x[18] , G3[17] , sum[18] ) ;
    _Psum _Psum_19( x[19] , G3[18] , sum[19] ) ;
    _Psum _Psum_20( x[20] , G3[19] , sum[20] ) ;
    _Psum _Psum_21( x[21] , G3[20] , sum[21] ) ;
    _Psum _Psum_22( x[22] , G3[21] , sum[22] ) ;
    _Psum _Psum_23( x[23] , G3[22] , sum[23] ) ;
    _Psum _Psum_24( x[24] , G3[23] , sum[24] ) ;
    _Psum _Psum_25( x[25] , G3[24] , sum[25] ) ;
    _Psum _Psum_26( x[26] , G3[25] , sum[26] ) ;
    _Psum _Psum_27( x[27] , G3[26] , sum[27] ) ;
    _Psum _Psum_28( x[28] , G3[27] , sum[28] ) ;
    _Psum _Psum_29( x[29] , G3[28] , sum[29] ) ;
    _Psum _Psum_30( x[30] , G3[29] , sum[30] ) ;
    _Psum _Psum_31( x[31] , G3[30] , sum[31] ) ;
    _Psum _Psum_32( x[32] , G3[31] , sum[32] ) ;
    _Psum _Psum_33( x[33] , G3[32] , sum[33] ) ;
    _Psum _Psum_34( x[34] , G3[33] , sum[34] ) ;
    _Psum _Psum_35( x[35] , G3[34] , sum[35] ) ;
    _Psum _Psum_36( x[36] , G3[35] , sum[36] ) ;
    _Psum _Psum_37( x[37] , G3[36] , sum[37] ) ;
    _Psum _Psum_38( x[38] , G3[37] , sum[38] ) ;
    _Psum _Psum_39( x[39] , G3[38] , sum[39] ) ;
    _Psum _Psum_40( x[40] , G3[39] , sum[40] ) ;
    _Psum _Psum_41( x[41] , G3[40] , sum[41] ) ;
    _Psum _Psum_42( x[42] , G3[41] , sum[42] ) ;
    _Psum _Psum_43( x[43] , G3[42] , sum[43] ) ;
    _Psum _Psum_44( x[44] , G3[43] , sum[44] ) ;
    _Psum _Psum_45( x[45] , G3[44] , sum[45] ) ;
    _Psum _Psum_46( x[46] , G3[45] , sum[46] ) ;
    _Psum _Psum_47( x[47] , G3[46] , sum[47] ) ;
    _Psum _Psum_48( x[48] , G3[47] , sum[48] ) ;
    _Psum _Psum_49( x[49] , G3[48] , sum[49] ) ;
    _Psum _Psum_50( x[50] , G3[49] , sum[50] ) ;
    _Psum _Psum_51( x[51] , G3[50] , sum[51] ) ;
    _Psum _Psum_52( x[52] , G3[51] , sum[52] ) ;
    _Psum _Psum_53( x[53] , G3[52] , sum[53] ) ;
    _Psum _Psum_54( x[54] , G3[53] , sum[54] ) ;
    _Psum _Psum_55( x[55] , G3[54] , sum[55] ) ;
    _Psum _Psum_56( x[56] , G3[55] , sum[56] ) ;
    _Psum _Psum_57( x[57] , G3[56] , sum[57] ) ;
    _Psum _Psum_58( x[58] , G3[57] , sum[58] ) ;
    _Psum _Psum_59( x[59] , G3[58] , sum[59] ) ;
    _Psum _Psum_60( x[60] , G3[59] , sum[60] ) ;
    _Psum _Psum_61( x[61] , G3[60] , sum[61] ) ;
    _Psum _Psum_62( x[62] , G3[61] , sum[62] ) ;
    _Psum _Psum_63( x[63] , G3[62] , sum[63] ) ;

endmodule
