module P32_node_adder(a, b, sum);
    input [31:0]a;
    input [31:0]b;
    output [31:0]sum;
    wire [31:0]g ;
    wire [31:0]p ;
    wire [31:0]x ;
    wire [31:0]G1 ;
    wire [31:0]G2 ;
    wire [31:0]G3 ;
    wire [31:0]Pr1 ;
    wire [31:0]Pr2 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;
    _gpx _gpx_16	(a[16],	b[16],	g[16], 	p[16], 	x[16]) ;
    _gpx _gpx_17	(a[17],	b[17],	g[17], 	p[17], 	x[17]) ;
    _gpx _gpx_18	(a[18],	b[18],	g[18], 	p[18], 	x[18]) ;
    _gpx _gpx_19	(a[19],	b[19],	g[19], 	p[19], 	x[19]) ;
    _gpx _gpx_20	(a[20],	b[20],	g[20], 	p[20], 	x[20]) ;
    _gpx _gpx_21	(a[21],	b[21],	g[21], 	p[21], 	x[21]) ;
    _gpx _gpx_22	(a[22],	b[22],	g[22], 	p[22], 	x[22]) ;
    _gpx _gpx_23	(a[23],	b[23],	g[23], 	p[23], 	x[23]) ;
    _gpx _gpx_24	(a[24],	b[24],	g[24], 	p[24], 	x[24]) ;
    _gpx _gpx_25	(a[25],	b[25],	g[25], 	p[25], 	x[25]) ;
    _gpx _gpx_26	(a[26],	b[26],	g[26], 	p[26], 	x[26]) ;
    _gpx _gpx_27	(a[27],	b[27],	g[27], 	p[27], 	x[27]) ;
    _gpx _gpx_28	(a[28],	b[28],	g[28], 	p[28], 	x[28]) ;
    _gpx _gpx_29	(a[29],	b[29],	g[29], 	p[29], 	x[29]) ;
    _gpx _gpx_30	(a[30],	b[30],	g[30], 	p[30], 	x[30]) ;
    _gpx _gpx_31	(a[31],	b[31],	g[31], 	p[31], 	x[31]) ;

    _2g1p_G2 _2g1p_G2_0( {g[0],g[31]} , p[0] , G1[0] ) ;
    _2g1p_G2 _2g1p_G2_1( {g[1],g[0]} , p[1] , G1[1] ) ;
    _2g1p_G2 _2g1p_G2_2( {g[2],g[1]} , p[2] , G1[2] ) ;
    _2g1p_G2 _2g1p_G2_3( {g[3],g[2]} , p[3] , G1[3] ) ;
    _2g1p_G2 _2g1p_G2_4( {g[4],g[3]} , p[4] , G1[4] ) ;
    _2g1p_G2 _2g1p_G2_5( {g[5],g[4]} , p[5] , G1[5] ) ;
    _2g1p_G2 _2g1p_G2_6( {g[6],g[5]} , p[6] , G1[6] ) ;
    _2g1p_G2 _2g1p_G2_7( {g[7],g[6]} , p[7] , G1[7] ) ;
    _2g1p_G2 _2g1p_G2_8( {g[8],g[7]} , p[8] , G1[8] ) ;
    _2g1p_G2 _2g1p_G2_9( {g[9],g[8]} , p[9] , G1[9] ) ;
    _2g1p_G2 _2g1p_G2_10( {g[10],g[9]} , p[10] , G1[10] ) ;
    _2g1p_G2 _2g1p_G2_11( {g[11],g[10]} , p[11] , G1[11] ) ;
    _2g1p_G2 _2g1p_G2_12( {g[12],g[11]} , p[12] , G1[12] ) ;
    _2g1p_G2 _2g1p_G2_13( {g[13],g[12]} , p[13] , G1[13] ) ;
    _2g1p_G2 _2g1p_G2_14( {g[14],g[13]} , p[14] , G1[14] ) ;
    _2g1p_G2 _2g1p_G2_15( {g[15],g[14]} , p[15] , G1[15] ) ;
    _2g1p_G2 _2g1p_G2_16( {g[16],g[15]} , p[16] , G1[16] ) ;
    _2g1p_G2 _2g1p_G2_17( {g[17],g[16]} , p[17] , G1[17] ) ;
    _2g1p_G2 _2g1p_G2_18( {g[18],g[17]} , p[18] , G1[18] ) ;
    _2g1p_G2 _2g1p_G2_19( {g[19],g[18]} , p[19] , G1[19] ) ;
    _2g1p_G2 _2g1p_G2_20( {g[20],g[19]} , p[20] , G1[20] ) ;
    _2g1p_G2 _2g1p_G2_21( {g[21],g[20]} , p[21] , G1[21] ) ;
    _2g1p_G2 _2g1p_G2_22( {g[22],g[21]} , p[22] , G1[22] ) ;
    _2g1p_G2 _2g1p_G2_23( {g[23],g[22]} , p[23] , G1[23] ) ;
    _2g1p_G2 _2g1p_G2_24( {g[24],g[23]} , p[24] , G1[24] ) ;
    _2g1p_G2 _2g1p_G2_25( {g[25],g[24]} , p[25] , G1[25] ) ;
    _2g1p_G2 _2g1p_G2_26( {g[26],g[25]} , p[26] , G1[26] ) ;
    _2g1p_G2 _2g1p_G2_27( {g[27],g[26]} , p[27] , G1[27] ) ;
    _2g1p_G2 _2g1p_G2_28( {g[28],g[27]} , p[28] , G1[28] ) ;
    _2g1p_G2 _2g1p_G2_29( {g[29],g[28]} , p[29] , G1[29] ) ;
    _2g1p_G2 _2g1p_G2_30( {g[30],g[29]} , p[30] , G1[30] ) ;
    _2g1p_G2 _2g1p_G2_31( {g[31],g[30]} , p[31] , G1[31] ) ;

    _2p_P2 _2p_P2_0( {p[0],p[31]} , Pr1[0] ) ;
    _2p_P2 _2p_P2_1( {p[1],p[0]} , Pr1[1] ) ;
    _2p_P2 _2p_P2_2( {p[2],p[1]} , Pr1[2] ) ;
    _2p_P2 _2p_P2_3( {p[3],p[2]} , Pr1[3] ) ;
    _2p_P2 _2p_P2_4( {p[4],p[3]} , Pr1[4] ) ;
    _2p_P2 _2p_P2_5( {p[5],p[4]} , Pr1[5] ) ;
    _2p_P2 _2p_P2_6( {p[6],p[5]} , Pr1[6] ) ;
    _2p_P2 _2p_P2_7( {p[7],p[6]} , Pr1[7] ) ;
    _2p_P2 _2p_P2_8( {p[8],p[7]} , Pr1[8] ) ;
    _2p_P2 _2p_P2_9( {p[9],p[8]} , Pr1[9] ) ;
    _2p_P2 _2p_P2_10( {p[10],p[9]} , Pr1[10] ) ;
    _2p_P2 _2p_P2_11( {p[11],p[10]} , Pr1[11] ) ;
    _2p_P2 _2p_P2_12( {p[12],p[11]} , Pr1[12] ) ;
    _2p_P2 _2p_P2_13( {p[13],p[12]} , Pr1[13] ) ;
    _2p_P2 _2p_P2_14( {p[14],p[13]} , Pr1[14] ) ;
    _2p_P2 _2p_P2_15( {p[15],p[14]} , Pr1[15] ) ;
    _2p_P2 _2p_P2_16( {p[16],p[15]} , Pr1[16] ) ;
    _2p_P2 _2p_P2_17( {p[17],p[16]} , Pr1[17] ) ;
    _2p_P2 _2p_P2_18( {p[18],p[17]} , Pr1[18] ) ;
    _2p_P2 _2p_P2_19( {p[19],p[18]} , Pr1[19] ) ;
    _2p_P2 _2p_P2_20( {p[20],p[19]} , Pr1[20] ) ;
    _2p_P2 _2p_P2_21( {p[21],p[20]} , Pr1[21] ) ;
    _2p_P2 _2p_P2_22( {p[22],p[21]} , Pr1[22] ) ;
    _2p_P2 _2p_P2_23( {p[23],p[22]} , Pr1[23] ) ;
    _2p_P2 _2p_P2_24( {p[24],p[23]} , Pr1[24] ) ;
    _2p_P2 _2p_P2_25( {p[25],p[24]} , Pr1[25] ) ;
    _2p_P2 _2p_P2_26( {p[26],p[25]} , Pr1[26] ) ;
    _2p_P2 _2p_P2_27( {p[27],p[26]} , Pr1[27] ) ;
    _2p_P2 _2p_P2_28( {p[28],p[27]} , Pr1[28] ) ;
    _2p_P2 _2p_P2_29( {p[29],p[28]} , Pr1[29] ) ;
    _2p_P2 _2p_P2_30( {p[30],p[29]} , Pr1[30] ) ;
    _2p_P2 _2p_P2_31( {p[31],p[30]} , Pr1[31] ) ;

    _4G3P_G4 _4G3P_G4_0( {G1[0],G1[30],G1[28],G1[26]} , {Pr1[0],Pr1[30],Pr1[28]} ,G2[0] ) ;
    _4G3P_G4 _4G3P_G4_1( {G1[1],G1[31],G1[29],G1[27]} , {Pr1[1],Pr1[31],Pr1[29]} ,G2[1] ) ;
    _4G3P_G4 _4G3P_G4_2( {G1[2],G1[0],G1[30],G1[28]} , {Pr1[2],Pr1[0],Pr1[30]} ,G2[2] ) ;
    _4G3P_G4 _4G3P_G4_3( {G1[3],G1[1],G1[31],G1[29]} , {Pr1[3],Pr1[1],Pr1[31]} ,G2[3] ) ;
    _4G3P_G4 _4G3P_G4_4( {G1[4],G1[2],G1[0],G1[30]} , {Pr1[4],Pr1[2],Pr1[0]} ,G2[4] ) ;
    _4G3P_G4 _4G3P_G4_5( {G1[5],G1[3],G1[1],G1[31]} , {Pr1[5],Pr1[3],Pr1[1]} ,G2[5] ) ;
    _4G3P_G4 _4G3P_G4_6( {G1[6],G1[4],G1[2],G1[0]} , {Pr1[6],Pr1[4],Pr1[2]} ,G2[6] ) ;
    _4G3P_G4 _4G3P_G4_7( {G1[7],G1[5],G1[3],G1[1]} , {Pr1[7],Pr1[5],Pr1[3]} ,G2[7] ) ;
    _4G3P_G4 _4G3P_G4_8( {G1[8],G1[6],G1[4],G1[2]} , {Pr1[8],Pr1[6],Pr1[4]} ,G2[8] ) ;
    _4G3P_G4 _4G3P_G4_9( {G1[9],G1[7],G1[5],G1[3]} , {Pr1[9],Pr1[7],Pr1[5]} ,G2[9] ) ;
    _4G3P_G4 _4G3P_G4_10( {G1[10],G1[8],G1[6],G1[4]} , {Pr1[10],Pr1[8],Pr1[6]} ,G2[10] ) ;
    _4G3P_G4 _4G3P_G4_11( {G1[11],G1[9],G1[7],G1[5]} , {Pr1[11],Pr1[9],Pr1[7]} ,G2[11] ) ;
    _4G3P_G4 _4G3P_G4_12( {G1[12],G1[10],G1[8],G1[6]} , {Pr1[12],Pr1[10],Pr1[8]} ,G2[12] ) ;
    _4G3P_G4 _4G3P_G4_13( {G1[13],G1[11],G1[9],G1[7]} , {Pr1[13],Pr1[11],Pr1[9]} ,G2[13] ) ;
    _4G3P_G4 _4G3P_G4_14( {G1[14],G1[12],G1[10],G1[8]} , {Pr1[14],Pr1[12],Pr1[10]} ,G2[14] ) ;
    _4G3P_G4 _4G3P_G4_15( {G1[15],G1[13],G1[11],G1[9]} , {Pr1[15],Pr1[13],Pr1[11]} ,G2[15] ) ;
    _4G3P_G4 _4G3P_G4_16( {G1[16],G1[14],G1[12],G1[10]} , {Pr1[16],Pr1[14],Pr1[12]} ,G2[16] ) ;
    _4G3P_G4 _4G3P_G4_17( {G1[17],G1[15],G1[13],G1[11]} , {Pr1[17],Pr1[15],Pr1[13]} ,G2[17] ) ;
    _4G3P_G4 _4G3P_G4_18( {G1[18],G1[16],G1[14],G1[12]} , {Pr1[18],Pr1[16],Pr1[14]} ,G2[18] ) ;
    _4G3P_G4 _4G3P_G4_19( {G1[19],G1[17],G1[15],G1[13]} , {Pr1[19],Pr1[17],Pr1[15]} ,G2[19] ) ;
    _4G3P_G4 _4G3P_G4_20( {G1[20],G1[18],G1[16],G1[14]} , {Pr1[20],Pr1[18],Pr1[16]} ,G2[20] ) ;
    _4G3P_G4 _4G3P_G4_21( {G1[21],G1[19],G1[17],G1[15]} , {Pr1[21],Pr1[19],Pr1[17]} ,G2[21] ) ;
    _4G3P_G4 _4G3P_G4_22( {G1[22],G1[20],G1[18],G1[16]} , {Pr1[22],Pr1[20],Pr1[18]} ,G2[22] ) ;
    _4G3P_G4 _4G3P_G4_23( {G1[23],G1[21],G1[19],G1[17]} , {Pr1[23],Pr1[21],Pr1[19]} ,G2[23] ) ;
    _4G3P_G4 _4G3P_G4_24( {G1[24],G1[22],G1[20],G1[18]} , {Pr1[24],Pr1[22],Pr1[20]} ,G2[24] ) ;
    _4G3P_G4 _4G3P_G4_25( {G1[25],G1[23],G1[21],G1[19]} , {Pr1[25],Pr1[23],Pr1[21]} ,G2[25] ) ;
    _4G3P_G4 _4G3P_G4_26( {G1[26],G1[24],G1[22],G1[20]} , {Pr1[26],Pr1[24],Pr1[22]} ,G2[26] ) ;
    _4G3P_G4 _4G3P_G4_27( {G1[27],G1[25],G1[23],G1[21]} , {Pr1[27],Pr1[25],Pr1[23]} ,G2[27] ) ;
    _4G3P_G4 _4G3P_G4_28( {G1[28],G1[26],G1[24],G1[22]} , {Pr1[28],Pr1[26],Pr1[24]} ,G2[28] ) ;
    _4G3P_G4 _4G3P_G4_29( {G1[29],G1[27],G1[25],G1[23]} , {Pr1[29],Pr1[27],Pr1[25]} ,G2[29] ) ;
    _4G3P_G4 _4G3P_G4_30( {G1[30],G1[28],G1[26],G1[24]} , {Pr1[30],Pr1[28],Pr1[26]} ,G2[30] ) ;
    _4G3P_G4 _4G3P_G4_31( {G1[31],G1[29],G1[27],G1[25]} , {Pr1[31],Pr1[29],Pr1[27]} ,G2[31] ) ;

    _P4 _P4_0( {Pr1[0],Pr1[30],Pr1[28],Pr1[26]} ,Pr2[0] ) ;
    _P4 _P4_1( {Pr1[1],Pr1[31],Pr1[29],Pr1[27]} ,Pr2[1] ) ;
    _P4 _P4_2( {Pr1[2],Pr1[0],Pr1[30],Pr1[28]} ,Pr2[2] ) ;
    _P4 _P4_3( {Pr1[3],Pr1[1],Pr1[31],Pr1[29]} ,Pr2[3] ) ;
    _P4 _P4_4( {Pr1[4],Pr1[2],Pr1[0],Pr1[30]} ,Pr2[4] ) ;
    _P4 _P4_5( {Pr1[5],Pr1[3],Pr1[1],Pr1[31]} ,Pr2[5] ) ;
    _P4 _P4_6( {Pr1[6],Pr1[4],Pr1[2],Pr1[0]} ,Pr2[6] ) ;
    _P4 _P4_7( {Pr1[7],Pr1[5],Pr1[3],Pr1[1]} ,Pr2[7] ) ;
    _P4 _P4_8( {Pr1[8],Pr1[6],Pr1[4],Pr1[2]} ,Pr2[8] ) ;
    _P4 _P4_9( {Pr1[9],Pr1[7],Pr1[5],Pr1[3]} ,Pr2[9] ) ;
    _P4 _P4_10( {Pr1[10],Pr1[8],Pr1[6],Pr1[4]} ,Pr2[10] ) ;
    _P4 _P4_11( {Pr1[11],Pr1[9],Pr1[7],Pr1[5]} ,Pr2[11] ) ;
    _P4 _P4_12( {Pr1[12],Pr1[10],Pr1[8],Pr1[6]} ,Pr2[12] ) ;
    _P4 _P4_13( {Pr1[13],Pr1[11],Pr1[9],Pr1[7]} ,Pr2[13] ) ;
    _P4 _P4_14( {Pr1[14],Pr1[12],Pr1[10],Pr1[8]} ,Pr2[14] ) ;
    _P4 _P4_15( {Pr1[15],Pr1[13],Pr1[11],Pr1[9]} ,Pr2[15] ) ;
    _P4 _P4_16( {Pr1[16],Pr1[14],Pr1[12],Pr1[10]} ,Pr2[16] ) ;
    _P4 _P4_17( {Pr1[17],Pr1[15],Pr1[13],Pr1[11]} ,Pr2[17] ) ;
    _P4 _P4_18( {Pr1[18],Pr1[16],Pr1[14],Pr1[12]} ,Pr2[18] ) ;
    _P4 _P4_19( {Pr1[19],Pr1[17],Pr1[15],Pr1[13]} ,Pr2[19] ) ;
    _P4 _P4_20( {Pr1[20],Pr1[18],Pr1[16],Pr1[14]} ,Pr2[20] ) ;
    _P4 _P4_21( {Pr1[21],Pr1[19],Pr1[17],Pr1[15]} ,Pr2[21] ) ;
    _P4 _P4_22( {Pr1[22],Pr1[20],Pr1[18],Pr1[16]} ,Pr2[22] ) ;
    _P4 _P4_23( {Pr1[23],Pr1[21],Pr1[19],Pr1[17]} ,Pr2[23] ) ;
    _P4 _P4_24( {Pr1[24],Pr1[22],Pr1[20],Pr1[18]} ,Pr2[24] ) ;
    _P4 _P4_25( {Pr1[25],Pr1[23],Pr1[21],Pr1[19]} ,Pr2[25] ) ;
    _P4 _P4_26( {Pr1[26],Pr1[24],Pr1[22],Pr1[20]} ,Pr2[26] ) ;
    _P4 _P4_27( {Pr1[27],Pr1[25],Pr1[23],Pr1[21]} ,Pr2[27] ) ;
    _P4 _P4_28( {Pr1[28],Pr1[26],Pr1[24],Pr1[22]} ,Pr2[28] ) ;
    _P4 _P4_29( {Pr1[29],Pr1[27],Pr1[25],Pr1[23]} ,Pr2[29] ) ;
    _P4 _P4_30( {Pr1[30],Pr1[28],Pr1[26],Pr1[24]} ,Pr2[30] ) ;
    _P4 _P4_31( {Pr1[31],Pr1[29],Pr1[27],Pr1[25]} ,Pr2[31] ) ;

    _4G3P_G4 _4G3P_G4_32( {G2[0],G2[24],G2[16],G2[8]} , {Pr2[0],Pr2[24],Pr2[16]} ,G3[0] ) ;
    _4G3P_G4 _4G3P_G4_33( {G2[1],G2[25],G2[17],G2[9]} , {Pr2[1],Pr2[25],Pr2[17]} ,G3[1] ) ;
    _4G3P_G4 _4G3P_G4_34( {G2[2],G2[26],G2[18],G2[10]} , {Pr2[2],Pr2[26],Pr2[18]} ,G3[2] ) ;
    _4G3P_G4 _4G3P_G4_35( {G2[3],G2[27],G2[19],G2[11]} , {Pr2[3],Pr2[27],Pr2[19]} ,G3[3] ) ;
    _4G3P_G4 _4G3P_G4_36( {G2[4],G2[28],G2[20],G2[12]} , {Pr2[4],Pr2[28],Pr2[20]} ,G3[4] ) ;
    _4G3P_G4 _4G3P_G4_37( {G2[5],G2[29],G2[21],G2[13]} , {Pr2[5],Pr2[29],Pr2[21]} ,G3[5] ) ;
    _4G3P_G4 _4G3P_G4_38( {G2[6],G2[30],G2[22],G2[14]} , {Pr2[6],Pr2[30],Pr2[22]} ,G3[6] ) ;
    _4G3P_G4 _4G3P_G4_39( {G2[7],G2[31],G2[23],G2[15]} , {Pr2[7],Pr2[31],Pr2[23]} ,G3[7] ) ;
    _4G3P_G4 _4G3P_G4_40( {G2[8],G2[0],G2[24],G2[16]} , {Pr2[8],Pr2[0],Pr2[24]} ,G3[8] ) ;
    _4G3P_G4 _4G3P_G4_41( {G2[9],G2[1],G2[25],G2[17]} , {Pr2[9],Pr2[1],Pr2[25]} ,G3[9] ) ;
    _4G3P_G4 _4G3P_G4_42( {G2[10],G2[2],G2[26],G2[18]} , {Pr2[10],Pr2[2],Pr2[26]} ,G3[10] ) ;
    _4G3P_G4 _4G3P_G4_43( {G2[11],G2[3],G2[27],G2[19]} , {Pr2[11],Pr2[3],Pr2[27]} ,G3[11] ) ;
    _4G3P_G4 _4G3P_G4_44( {G2[12],G2[4],G2[28],G2[20]} , {Pr2[12],Pr2[4],Pr2[28]} ,G3[12] ) ;
    _4G3P_G4 _4G3P_G4_45( {G2[13],G2[5],G2[29],G2[21]} , {Pr2[13],Pr2[5],Pr2[29]} ,G3[13] ) ;
    _4G3P_G4 _4G3P_G4_46( {G2[14],G2[6],G2[30],G2[22]} , {Pr2[14],Pr2[6],Pr2[30]} ,G3[14] ) ;
    _4G3P_G4 _4G3P_G4_47( {G2[15],G2[7],G2[31],G2[23]} , {Pr2[15],Pr2[7],Pr2[31]} ,G3[15] ) ;
    _4G3P_G4 _4G3P_G4_48( {G2[16],G2[8],G2[0],G2[24]} , {Pr2[16],Pr2[8],Pr2[0]} ,G3[16] ) ;
    _4G3P_G4 _4G3P_G4_49( {G2[17],G2[9],G2[1],G2[25]} , {Pr2[17],Pr2[9],Pr2[1]} ,G3[17] ) ;
    _4G3P_G4 _4G3P_G4_50( {G2[18],G2[10],G2[2],G2[26]} , {Pr2[18],Pr2[10],Pr2[2]} ,G3[18] ) ;
    _4G3P_G4 _4G3P_G4_51( {G2[19],G2[11],G2[3],G2[27]} , {Pr2[19],Pr2[11],Pr2[3]} ,G3[19] ) ;
    _4G3P_G4 _4G3P_G4_52( {G2[20],G2[12],G2[4],G2[28]} , {Pr2[20],Pr2[12],Pr2[4]} ,G3[20] ) ;
    _4G3P_G4 _4G3P_G4_53( {G2[21],G2[13],G2[5],G2[29]} , {Pr2[21],Pr2[13],Pr2[5]} ,G3[21] ) ;
    _4G3P_G4 _4G3P_G4_54( {G2[22],G2[14],G2[6],G2[30]} , {Pr2[22],Pr2[14],Pr2[6]} ,G3[22] ) ;
    _4G3P_G4 _4G3P_G4_55( {G2[23],G2[15],G2[7],G2[31]} , {Pr2[23],Pr2[15],Pr2[7]} ,G3[23] ) ;
    _4G3P_G4 _4G3P_G4_56( {G2[24],G2[16],G2[8],G2[0]} , {Pr2[24],Pr2[16],Pr2[8]} ,G3[24] ) ;
    _4G3P_G4 _4G3P_G4_57( {G2[25],G2[17],G2[9],G2[1]} , {Pr2[25],Pr2[17],Pr2[9]} ,G3[25] ) ;
    _4G3P_G4 _4G3P_G4_58( {G2[26],G2[18],G2[10],G2[2]} , {Pr2[26],Pr2[18],Pr2[10]} ,G3[26] ) ;
    _4G3P_G4 _4G3P_G4_59( {G2[27],G2[19],G2[11],G2[3]} , {Pr2[27],Pr2[19],Pr2[11]} ,G3[27] ) ;
    _4G3P_G4 _4G3P_G4_60( {G2[28],G2[20],G2[12],G2[4]} , {Pr2[28],Pr2[20],Pr2[12]} ,G3[28] ) ;
    _4G3P_G4 _4G3P_G4_61( {G2[29],G2[21],G2[13],G2[5]} , {Pr2[29],Pr2[21],Pr2[13]} ,G3[29] ) ;
    _4G3P_G4 _4G3P_G4_62( {G2[30],G2[22],G2[14],G2[6]} , {Pr2[30],Pr2[22],Pr2[14]} ,G3[30] ) ;
    _4G3P_G4 _4G3P_G4_63( {G2[31],G2[23],G2[15],G2[7]} , {Pr2[31],Pr2[23],Pr2[15]} ,G3[31] ) ;

    _Psum _Psum_0( x[0] , G3[31] , sum[0] ) ;
    _Psum _Psum_1( x[1] , G3[0] , sum[1] ) ;
    _Psum _Psum_2( x[2] , G3[1] , sum[2] ) ;
    _Psum _Psum_3( x[3] , G3[2] , sum[3] ) ;
    _Psum _Psum_4( x[4] , G3[3] , sum[4] ) ;
    _Psum _Psum_5( x[5] , G3[4] , sum[5] ) ;
    _Psum _Psum_6( x[6] , G3[5] , sum[6] ) ;
    _Psum _Psum_7( x[7] , G3[6] , sum[7] ) ;
    _Psum _Psum_8( x[8] , G3[7] , sum[8] ) ;
    _Psum _Psum_9( x[9] , G3[8] , sum[9] ) ;
    _Psum _Psum_10( x[10] , G3[9] , sum[10] ) ;
    _Psum _Psum_11( x[11] , G3[10] , sum[11] ) ;
    _Psum _Psum_12( x[12] , G3[11] , sum[12] ) ;
    _Psum _Psum_13( x[13] , G3[12] , sum[13] ) ;
    _Psum _Psum_14( x[14] , G3[13] , sum[14] ) ;
    _Psum _Psum_15( x[15] , G3[14] , sum[15] ) ;
    _Psum _Psum_16( x[16] , G3[15] , sum[16] ) ;
    _Psum _Psum_17( x[17] , G3[16] , sum[17] ) ;
    _Psum _Psum_18( x[18] , G3[17] , sum[18] ) ;
    _Psum _Psum_19( x[19] , G3[18] , sum[19] ) ;
    _Psum _Psum_20( x[20] , G3[19] , sum[20] ) ;
    _Psum _Psum_21( x[21] , G3[20] , sum[21] ) ;
    _Psum _Psum_22( x[22] , G3[21] , sum[22] ) ;
    _Psum _Psum_23( x[23] , G3[22] , sum[23] ) ;
    _Psum _Psum_24( x[24] , G3[23] , sum[24] ) ;
    _Psum _Psum_25( x[25] , G3[24] , sum[25] ) ;
    _Psum _Psum_26( x[26] , G3[25] , sum[26] ) ;
    _Psum _Psum_27( x[27] , G3[26] , sum[27] ) ;
    _Psum _Psum_28( x[28] , G3[27] , sum[28] ) ;
    _Psum _Psum_29( x[29] , G3[28] , sum[29] ) ;
    _Psum _Psum_30( x[30] , G3[29] , sum[30] ) ;
    _Psum _Psum_31( x[31] , G3[30] , sum[31] ) ;

endmodule
