// 1. _gpx(a, b, g, p, x)
// 2. _4g2p_R4(g, p, R)
// 3. _4p_Q4((p, Q)
// 4. _4R2Q_R4(R_in, Q_in, R_out)
// 5. _D16(R, p, D)
// 6. _Jsum(R, D, x, sum)
// 7. _1R4Q_Q4(R_in, Q_in, Q_out)
// 8. _D64_1(p, g, D)
// 9. _D64_2(D_in, R_in, Q_in, D_out)
// 10._2g_R2(g,R)
// 11._2p_Q2(p,Q)
// 12._4g2p_H4(g, p, H)
// 13._P4(p_in,p_out)
// 14._4G3P_G4(G_in, P_in, G_out)
// 15._Lsum(p, x, H, sum)
// 16._2g_H2(g, H)
// 17._2p_P2(p, Pr)
// 18._Psum(x, G, sum)
// 19._2g1p_G2(g, p, G_out)
// 20._2R1Q_R2(R_in, Q_in, R_out)
// 21._Psum_sparse2(x, g, p, G, sum)
// 22._Lsum_sparse2(x, g, p, H, sum)
// 23._Jsum_sparse2(g, p, R ,D , x, sum )


// .1
//-------------------------------------------------------
module _gpx(a, b, g, p, x);

    input a;
    input b;
    output g;
    output p;
    output x;
    
    assign p = a | b ;
    assign g = a & b ;
    assign x = a ^ b ;

endmodule



// .2
//-------------------------------------------------------
module _4g2p_R4(g, p, R);

    input [3:0]g;
    input [1:0]p;
    output R;
    
    assign R =  g[3] |
                g[2] |
                p[1] & g[1] |
                p[1] & p[0] & g[0] ;
endmodule



// .3
//-------------------------------------------------------
module _4p_Q4(p, Q);

    input [3:0]p;
    output Q;
    
    assign Q = p[3] & p[2] & p[1] & p[0];
    
endmodule



// .4
//-------------------------------------------------------
module _4R2Q_R4(R_in, Q_in, R_out);

    input [3:0]R_in;
    input [1:0]Q_in;
    output R_out;
    
    assign  R_out = R_in[3] |
                    R_in[2] |
                    Q_in[1] & R_in[1] |
                    Q_in[1] & Q_in[0] & R_in[0] ;

endmodule



// .5
//-------------------------------------------------------
module _D16(p, R, Q, D);


    input [1:0]p;
    input R;
    input Q;
    output D;
    
    assign D = (p[1] & R) | (p[0] & Q) ;

endmodule



// .6
//-------------------------------------------------------
module _Jsum(R, D, x, sum);

    input R;
    input D;
    input x;
    output sum;

    assign sum = R ? (x ^ D) : x ;
    
endmodule



// .7
//-------------------------------------------------------
module _1R4Q_Q4(R_in, Q_in, Q_out);

    input R_in;
    input [3:0]Q_in;
    output Q_out;
    
    assign Q_out =  Q_in[3] &
                    Q_in[2] &
                    Q_in[1] &
                    ( Q_in[0] | R_in ) ;
endmodule



// .8
//-------------------------------------------------------
module _D64_1(p, g, D);
    
    input [2:0]p;
    input [1:0]g;
    output D ;
    
    assign D =  g[1] |
                g[0] & p[2] |
                p[2] & p[1] & p[0] ;

endmodule



// .9
//-------------------------------------------------------
module _D64_2(D_in, R_in, Q_in, D_out);
    
    input D_in;
    input R_in;
    input Q_in;
    output D_out;
    
    assign D_out = D_in & ( R_in | Q_in ) ;

endmodule



// .10
//-------------------------------------------------------
module _2g_R2(g,R);
    
    input [1:0]g;
    output R;
    
    assign R = g[1] | g[0] ;
    
endmodule



// .11
//-------------------------------------------------------
module _2p_Q2(p,Q);
    
    input [1:0]p;
    output Q;
    
    assign Q = p[1] & p[0] ;
    
endmodule



// .12
//-------------------------------------------------------
module _4g2p_H4(g, p, H);

    input [3:0]g;
    input [1:0]p;
    output H;
    
    assign H = g[3] | g[2] | p[1]&g[1] | p[1]&p[0]&g[0] ;

endmodule



// .13
//-------------------------------------------------------
module _P4(p_in,p_out);

    input [3:0]p_in;
    output p_out;
    
    assign p_out = p_in[3] & p_in[2] & p_in[1] & p_in[0] ;
    
endmodule



// .14
//-------------------------------------------------------
module _4G3P_G4(G_in, P_in, G_out);

    input [3:0]G_in;
    input [2:0]P_in;
    output G_out;
    
    assign G_out =  G_in[3] | 
                    P_in[2] & G_in[2] | 
                    P_in[2] & P_in[1] & G_in[1] | 
                    P_in[2] & P_in[1] & P_in[0] & G_in[0];

endmodule



// .15
//-------------------------------------------------------
module _Lsum(p, x, H, sum);

    input p;
    input x;
    input H;
    output sum;

    assign sum = H ? (x ^ p) : x ;
    
endmodule



// .16
//-------------------------------------------------------
module _2g_H2(g, H);

    input [1:0]g;
    output H;
    
    assign H = g[1] | g[0] ;

endmodule



// .17
//-------------------------------------------------------
module _2p_P2(p, Pr);

    input [1:0]p;
    output Pr;
    
    assign Pr = p[1] & p[0] ;

endmodule




// .18
//-------------------------------------------------------
module _Psum(x, G, sum);

    input x;
    input G;
    output sum;

    assign sum = G ^ x ;
    
endmodule



// .19
//-------------------------------------------------------
module _2g1p_G2(g, p, G_out);
    
    input [1:0]g;
    input p;
    output G_out;

    assign G_out = g[1] | p & g[0] ;
endmodule



// .20
//-------------------------------------------------------
module _2R1Q_R2(R_in, Q_in, R_out);
    
    input [1:0]R_in;
    input Q_in;
    output R_out;
    
    assign R_out = R_in[1] | Q_in & R_in[0] ;

endmodule



// .21
//-------------------------------------------------------
module _Psum_sparse2(x, g, p, G, sum);
    
    input [1:0]x;
    input g;
    input p;
    input G;
    output [1:0]sum;

    assign sum[0] = G ^ x[0] ;
    assign sum[1] = x[1] ^ ( g | (p & G) ) ;
    
endmodule



// .22
//-------------------------------------------------------
module _Lsum_sparse2(x, g, p, H, sum);
    
    input [1:0]x;
    input g;
    input [1:0]p;
    input H;
    output [1:0]sum;

    assign sum[0] = H ? (x[0] ^ p[0]) : x[0] ;
    assign sum[1] = H ? (x[1] ^ (g | p[1] & p[0])) : (x[1] ^ g) ;
    
endmodule




// .23
//-------------------------------------------------------
module _Jsum_sparse2(g, p, R ,D , x, sum );
    
    input g;
    input p;
    input R;
    input D;
    input [1:0]x;    
    output [1:0]sum;
    
    assign sum[0] = R ? (x[0] ^ D) : x[0] ;
    assign sum[1] = R ? (x[1] ^ (g | p&D)) : x[1]^g ;
    
endmodule




// .24
//-------------------------------------------------------
module _Psum_sparse4(x, g, p, G, sum);
    
    input [3:0]x;
    input [2:0]g;
    input [2:0]p;
    input G;
    output [3:0]sum;

    assign sum[0] = G ^ x[0] ;
    assign sum[1] = x[1] ^ ( g[0] | (p[0] & G) ) ;
    assign sum[2] = x[2] ^ ( g[1] | (p[1] & g[0]) | (p[1]&p[0]&G)) ;
    assign sum[3] = x[3] ^ ( g[2] | (p[2] & g[1]) | ( p[2] & p[1] & g[0]) | (p[2]&p[1]&p[0]&G)) ;
    
endmodule




// .25
//-------------------------------------------------------
module _Lsum_sparse4(x, g, p, H, sum);
    
    input [3:0]x;
    input [2:0]g;
    input [3:0]p;
    input H;
    output [3:0]sum;

    assign sum[0] = H ? (x[0] ^ p[0]) : x[0] ;
    assign sum[1] = H ? (x[1] ^ (g[0] | (p[1]&p[0]) )) : (x[1] ^ g[0]) ;
    assign sum[2] = H ? (x[2] ^ (g[1] | (p[2]&g[0]) | (p[2]&p[1]&p[0]) )) : (x[2] ^ (g[1] | (p[2]&g[0])) ) ;
    assign sum[3] = H ? (x[3] ^ (g[2] | (p[3]&g[1]) | (p[3]&p[2]&g[0]) | (p[3]&p[2]&p[1]&p[0]) )) : (x[3] ^ (g[2] | (p[3]&g[1]) | (p[3]&p[2]&g[0]) )) ;
endmodule



// .26
//-------------------------------------------------------
module _Jsum_sparse4(g, p, R ,D , x, sum );
    
    input [2:0]g;
    input [2:0]p;
    input R;
    input D;
    input [3:0]x;    
    output [3:0]sum;
    
    assign sum[0] = R ? (x[0] ^ D) : x[0] ;
    assign sum[1] = R ? (x[1] ^ (g[0] | p[0]&D)) : x[1]^g[0] ;
    assign sum[2] = R ? (x[2] ^ (g[1] | p[1]&g[0] | p[1]&p[0]&D)) : x[2] ^ (g[1] | p[1]&g[0]) ;
    assign sum[3] = R ? (x[3] ^ (g[2] | p[2]&g[1] | p[2]&p[1]&g[0] | p[2]&p[1]&p[0]&D)) : x[3] ^ ( g[2] | p[2]&g[1] | p[2]&p[1]&g[0] ) ;

endmodule






