module J64_node_adder(a, b, sum);
    input [63:0]a;
    input [63:0]b;
    output [63:0]sum;
    wire [63:0]g ;
    wire [63:0]p ;
    wire [63:0]x ;
    wire [63:0]R1 ;
    wire [63:0]R2 ;
    wire [63:0]R3 ;
    wire [63:0]Q1 ;
    wire [63:0]Q2 ;
    wire [63:0]D1 ;
    wire [63:0]D2 ;
    wire [63:0]D3 ;

    _gpx _gpx_0	(a[0],	b[0],	g[0], 	p[0], 	x[0]) ;
    _gpx _gpx_1	(a[1],	b[1],	g[1], 	p[1], 	x[1]) ;
    _gpx _gpx_2	(a[2],	b[2],	g[2], 	p[2], 	x[2]) ;
    _gpx _gpx_3	(a[3],	b[3],	g[3], 	p[3], 	x[3]) ;
    _gpx _gpx_4	(a[4],	b[4],	g[4], 	p[4], 	x[4]) ;
    _gpx _gpx_5	(a[5],	b[5],	g[5], 	p[5], 	x[5]) ;
    _gpx _gpx_6	(a[6],	b[6],	g[6], 	p[6], 	x[6]) ;
    _gpx _gpx_7	(a[7],	b[7],	g[7], 	p[7], 	x[7]) ;
    _gpx _gpx_8	(a[8],	b[8],	g[8], 	p[8], 	x[8]) ;
    _gpx _gpx_9	(a[9],	b[9],	g[9], 	p[9], 	x[9]) ;
    _gpx _gpx_10	(a[10],	b[10],	g[10], 	p[10], 	x[10]) ;
    _gpx _gpx_11	(a[11],	b[11],	g[11], 	p[11], 	x[11]) ;
    _gpx _gpx_12	(a[12],	b[12],	g[12], 	p[12], 	x[12]) ;
    _gpx _gpx_13	(a[13],	b[13],	g[13], 	p[13], 	x[13]) ;
    _gpx _gpx_14	(a[14],	b[14],	g[14], 	p[14], 	x[14]) ;
    _gpx _gpx_15	(a[15],	b[15],	g[15], 	p[15], 	x[15]) ;
    _gpx _gpx_16	(a[16],	b[16],	g[16], 	p[16], 	x[16]) ;
    _gpx _gpx_17	(a[17],	b[17],	g[17], 	p[17], 	x[17]) ;
    _gpx _gpx_18	(a[18],	b[18],	g[18], 	p[18], 	x[18]) ;
    _gpx _gpx_19	(a[19],	b[19],	g[19], 	p[19], 	x[19]) ;
    _gpx _gpx_20	(a[20],	b[20],	g[20], 	p[20], 	x[20]) ;
    _gpx _gpx_21	(a[21],	b[21],	g[21], 	p[21], 	x[21]) ;
    _gpx _gpx_22	(a[22],	b[22],	g[22], 	p[22], 	x[22]) ;
    _gpx _gpx_23	(a[23],	b[23],	g[23], 	p[23], 	x[23]) ;
    _gpx _gpx_24	(a[24],	b[24],	g[24], 	p[24], 	x[24]) ;
    _gpx _gpx_25	(a[25],	b[25],	g[25], 	p[25], 	x[25]) ;
    _gpx _gpx_26	(a[26],	b[26],	g[26], 	p[26], 	x[26]) ;
    _gpx _gpx_27	(a[27],	b[27],	g[27], 	p[27], 	x[27]) ;
    _gpx _gpx_28	(a[28],	b[28],	g[28], 	p[28], 	x[28]) ;
    _gpx _gpx_29	(a[29],	b[29],	g[29], 	p[29], 	x[29]) ;
    _gpx _gpx_30	(a[30],	b[30],	g[30], 	p[30], 	x[30]) ;
    _gpx _gpx_31	(a[31],	b[31],	g[31], 	p[31], 	x[31]) ;
    _gpx _gpx_32	(a[32],	b[32],	g[32], 	p[32], 	x[32]) ;
    _gpx _gpx_33	(a[33],	b[33],	g[33], 	p[33], 	x[33]) ;
    _gpx _gpx_34	(a[34],	b[34],	g[34], 	p[34], 	x[34]) ;
    _gpx _gpx_35	(a[35],	b[35],	g[35], 	p[35], 	x[35]) ;
    _gpx _gpx_36	(a[36],	b[36],	g[36], 	p[36], 	x[36]) ;
    _gpx _gpx_37	(a[37],	b[37],	g[37], 	p[37], 	x[37]) ;
    _gpx _gpx_38	(a[38],	b[38],	g[38], 	p[38], 	x[38]) ;
    _gpx _gpx_39	(a[39],	b[39],	g[39], 	p[39], 	x[39]) ;
    _gpx _gpx_40	(a[40],	b[40],	g[40], 	p[40], 	x[40]) ;
    _gpx _gpx_41	(a[41],	b[41],	g[41], 	p[41], 	x[41]) ;
    _gpx _gpx_42	(a[42],	b[42],	g[42], 	p[42], 	x[42]) ;
    _gpx _gpx_43	(a[43],	b[43],	g[43], 	p[43], 	x[43]) ;
    _gpx _gpx_44	(a[44],	b[44],	g[44], 	p[44], 	x[44]) ;
    _gpx _gpx_45	(a[45],	b[45],	g[45], 	p[45], 	x[45]) ;
    _gpx _gpx_46	(a[46],	b[46],	g[46], 	p[46], 	x[46]) ;
    _gpx _gpx_47	(a[47],	b[47],	g[47], 	p[47], 	x[47]) ;
    _gpx _gpx_48	(a[48],	b[48],	g[48], 	p[48], 	x[48]) ;
    _gpx _gpx_49	(a[49],	b[49],	g[49], 	p[49], 	x[49]) ;
    _gpx _gpx_50	(a[50],	b[50],	g[50], 	p[50], 	x[50]) ;
    _gpx _gpx_51	(a[51],	b[51],	g[51], 	p[51], 	x[51]) ;
    _gpx _gpx_52	(a[52],	b[52],	g[52], 	p[52], 	x[52]) ;
    _gpx _gpx_53	(a[53],	b[53],	g[53], 	p[53], 	x[53]) ;
    _gpx _gpx_54	(a[54],	b[54],	g[54], 	p[54], 	x[54]) ;
    _gpx _gpx_55	(a[55],	b[55],	g[55], 	p[55], 	x[55]) ;
    _gpx _gpx_56	(a[56],	b[56],	g[56], 	p[56], 	x[56]) ;
    _gpx _gpx_57	(a[57],	b[57],	g[57], 	p[57], 	x[57]) ;
    _gpx _gpx_58	(a[58],	b[58],	g[58], 	p[58], 	x[58]) ;
    _gpx _gpx_59	(a[59],	b[59],	g[59], 	p[59], 	x[59]) ;
    _gpx _gpx_60	(a[60],	b[60],	g[60], 	p[60], 	x[60]) ;
    _gpx _gpx_61	(a[61],	b[61],	g[61], 	p[61], 	x[61]) ;
    _gpx _gpx_62	(a[62],	b[62],	g[62], 	p[62], 	x[62]) ;
    _gpx _gpx_63	(a[63],	b[63],	g[63], 	p[63], 	x[63]) ;

    _4g2p_R4 _4g2p_R4_1	( {g[1],g[0],g[63],g[62]} ,	{p[0],p[63]} ,	R1[1] ) ;
    _4g2p_R4 _4g2p_R4_3	( {g[3],g[2],g[1],g[0]} ,	{p[2],p[1]} ,	R1[3] ) ;
    _4g2p_R4 _4g2p_R4_5	( {g[5],g[4],g[3],g[2]} ,	{p[4],p[3]} ,	R1[5] ) ;
    _4g2p_R4 _4g2p_R4_7	( {g[7],g[6],g[5],g[4]} ,	{p[6],p[5]} ,	R1[7] ) ;
    _4g2p_R4 _4g2p_R4_9	( {g[9],g[8],g[7],g[6]} ,	{p[8],p[7]} ,	R1[9] ) ;
    _4g2p_R4 _4g2p_R4_11	( {g[11],g[10],g[9],g[8]} ,	{p[10],p[9]} ,	R1[11] ) ;
    _4g2p_R4 _4g2p_R4_13	( {g[13],g[12],g[11],g[10]} ,	{p[12],p[11]} ,	R1[13] ) ;
    _4g2p_R4 _4g2p_R4_15	( {g[15],g[14],g[13],g[12]} ,	{p[14],p[13]} ,	R1[15] ) ;
    _4g2p_R4 _4g2p_R4_17	( {g[17],g[16],g[15],g[14]} ,	{p[16],p[15]} ,	R1[17] ) ;
    _4g2p_R4 _4g2p_R4_19	( {g[19],g[18],g[17],g[16]} ,	{p[18],p[17]} ,	R1[19] ) ;
    _4g2p_R4 _4g2p_R4_21	( {g[21],g[20],g[19],g[18]} ,	{p[20],p[19]} ,	R1[21] ) ;
    _4g2p_R4 _4g2p_R4_23	( {g[23],g[22],g[21],g[20]} ,	{p[22],p[21]} ,	R1[23] ) ;
    _4g2p_R4 _4g2p_R4_25	( {g[25],g[24],g[23],g[22]} ,	{p[24],p[23]} ,	R1[25] ) ;
    _4g2p_R4 _4g2p_R4_27	( {g[27],g[26],g[25],g[24]} ,	{p[26],p[25]} ,	R1[27] ) ;
    _4g2p_R4 _4g2p_R4_29	( {g[29],g[28],g[27],g[26]} ,	{p[28],p[27]} ,	R1[29] ) ;
    _4g2p_R4 _4g2p_R4_31	( {g[31],g[30],g[29],g[28]} ,	{p[30],p[29]} ,	R1[31] ) ;
    _4g2p_R4 _4g2p_R4_33	( {g[33],g[32],g[31],g[30]} ,	{p[32],p[31]} ,	R1[33] ) ;
    _4g2p_R4 _4g2p_R4_35	( {g[35],g[34],g[33],g[32]} ,	{p[34],p[33]} ,	R1[35] ) ;
    _4g2p_R4 _4g2p_R4_37	( {g[37],g[36],g[35],g[34]} ,	{p[36],p[35]} ,	R1[37] ) ;
    _4g2p_R4 _4g2p_R4_39	( {g[39],g[38],g[37],g[36]} ,	{p[38],p[37]} ,	R1[39] ) ;
    _4g2p_R4 _4g2p_R4_41	( {g[41],g[40],g[39],g[38]} ,	{p[40],p[39]} ,	R1[41] ) ;
    _4g2p_R4 _4g2p_R4_43	( {g[43],g[42],g[41],g[40]} ,	{p[42],p[41]} ,	R1[43] ) ;
    _4g2p_R4 _4g2p_R4_45	( {g[45],g[44],g[43],g[42]} ,	{p[44],p[43]} ,	R1[45] ) ;
    _4g2p_R4 _4g2p_R4_47	( {g[47],g[46],g[45],g[44]} ,	{p[46],p[45]} ,	R1[47] ) ;
    _4g2p_R4 _4g2p_R4_49	( {g[49],g[48],g[47],g[46]} ,	{p[48],p[47]} ,	R1[49] ) ;
    _4g2p_R4 _4g2p_R4_51	( {g[51],g[50],g[49],g[48]} ,	{p[50],p[49]} ,	R1[51] ) ;
    _4g2p_R4 _4g2p_R4_53	( {g[53],g[52],g[51],g[50]} ,	{p[52],p[51]} ,	R1[53] ) ;
    _4g2p_R4 _4g2p_R4_55	( {g[55],g[54],g[53],g[52]} ,	{p[54],p[53]} ,	R1[55] ) ;
    _4g2p_R4 _4g2p_R4_57	( {g[57],g[56],g[55],g[54]} ,	{p[56],p[55]} ,	R1[57] ) ;
    _4g2p_R4 _4g2p_R4_59	( {g[59],g[58],g[57],g[56]} ,	{p[58],p[57]} ,	R1[59] ) ;
    _4g2p_R4 _4g2p_R4_61	( {g[61],g[60],g[59],g[58]} ,	{p[60],p[59]} ,	R1[61] ) ;
    _4g2p_R4 _4g2p_R4_63	( {g[63],g[62],g[61],g[60]} ,	{p[62],p[61]} ,	R1[63] ) ;

    _4p_Q4 _4p_Q4_0	({p[0],	p[63],	p[62],	p[61]} ,	Q1[0] ) ;
    _4p_Q4 _4p_Q4_2	({p[2],	p[1],	p[0],	p[63]} ,	Q1[2] ) ;
    _4p_Q4 _4p_Q4_4	({p[4],	p[3],	p[2],	p[1]} ,	Q1[4] ) ;
    _4p_Q4 _4p_Q4_6	({p[6],	p[5],	p[4],	p[3]} ,	Q1[6] ) ;
    _4p_Q4 _4p_Q4_8	({p[8],	p[7],	p[6],	p[5]} ,	Q1[8] ) ;
    _4p_Q4 _4p_Q4_10	({p[10],	p[9],	p[8],	p[7]} ,	Q1[10] ) ;
    _4p_Q4 _4p_Q4_12	({p[12],	p[11],	p[10],	p[9]} ,	Q1[12] ) ;
    _4p_Q4 _4p_Q4_14	({p[14],	p[13],	p[12],	p[11]} ,	Q1[14] ) ;
    _4p_Q4 _4p_Q4_16	({p[16],	p[15],	p[14],	p[13]} ,	Q1[16] ) ;
    _4p_Q4 _4p_Q4_18	({p[18],	p[17],	p[16],	p[15]} ,	Q1[18] ) ;
    _4p_Q4 _4p_Q4_20	({p[20],	p[19],	p[18],	p[17]} ,	Q1[20] ) ;
    _4p_Q4 _4p_Q4_22	({p[22],	p[21],	p[20],	p[19]} ,	Q1[22] ) ;
    _4p_Q4 _4p_Q4_24	({p[24],	p[23],	p[22],	p[21]} ,	Q1[24] ) ;
    _4p_Q4 _4p_Q4_26	({p[26],	p[25],	p[24],	p[23]} ,	Q1[26] ) ;
    _4p_Q4 _4p_Q4_28	({p[28],	p[27],	p[26],	p[25]} ,	Q1[28] ) ;
    _4p_Q4 _4p_Q4_30	({p[30],	p[29],	p[28],	p[27]} ,	Q1[30] ) ;
    _4p_Q4 _4p_Q4_32	({p[32],	p[31],	p[30],	p[29]} ,	Q1[32] ) ;
    _4p_Q4 _4p_Q4_34	({p[34],	p[33],	p[32],	p[31]} ,	Q1[34] ) ;
    _4p_Q4 _4p_Q4_36	({p[36],	p[35],	p[34],	p[33]} ,	Q1[36] ) ;
    _4p_Q4 _4p_Q4_38	({p[38],	p[37],	p[36],	p[35]} ,	Q1[38] ) ;
    _4p_Q4 _4p_Q4_40	({p[40],	p[39],	p[38],	p[37]} ,	Q1[40] ) ;
    _4p_Q4 _4p_Q4_42	({p[42],	p[41],	p[40],	p[39]} ,	Q1[42] ) ;
    _4p_Q4 _4p_Q4_44	({p[44],	p[43],	p[42],	p[41]} ,	Q1[44] ) ;
    _4p_Q4 _4p_Q4_46	({p[46],	p[45],	p[44],	p[43]} ,	Q1[46] ) ;
    _4p_Q4 _4p_Q4_48	({p[48],	p[47],	p[46],	p[45]} ,	Q1[48] ) ;
    _4p_Q4 _4p_Q4_50	({p[50],	p[49],	p[48],	p[47]} ,	Q1[50] ) ;
    _4p_Q4 _4p_Q4_52	({p[52],	p[51],	p[50],	p[49]} ,	Q1[52] ) ;
    _4p_Q4 _4p_Q4_54	({p[54],	p[53],	p[52],	p[51]} ,	Q1[54] ) ;
    _4p_Q4 _4p_Q4_56	({p[56],	p[55],	p[54],	p[53]} ,	Q1[56] ) ;
    _4p_Q4 _4p_Q4_58	({p[58],	p[57],	p[56],	p[55]} ,	Q1[58] ) ;
    _4p_Q4 _4p_Q4_60	({p[60],	p[59],	p[58],	p[57]} ,	Q1[60] ) ;
    _4p_Q4 _4p_Q4_62	({p[62],	p[61],	p[60],	p[59]} ,	Q1[62] ) ;

    _4R2Q_R4 _4R2Q_R4_1( {R1[1],R1[61],R1[57],R1[53] }, {Q1[60],Q1[56]} ,R2[1] ) ;
    _4R2Q_R4 _4R2Q_R4_3( {R1[3],R1[63],R1[59],R1[55] }, {Q1[62],Q1[58]} ,R2[3] ) ;
    _4R2Q_R4 _4R2Q_R4_5( {R1[5],R1[1],R1[61],R1[57] }, {Q1[0],Q1[60]} ,R2[5] ) ;
    _4R2Q_R4 _4R2Q_R4_7( {R1[7],R1[3],R1[63],R1[59] }, {Q1[2],Q1[62]} ,R2[7] ) ;
    _4R2Q_R4 _4R2Q_R4_9( {R1[9],R1[5],R1[1],R1[61] }, {Q1[4],Q1[0]} ,R2[9] ) ;
    _4R2Q_R4 _4R2Q_R4_11( {R1[11],R1[7],R1[3],R1[63] }, {Q1[6],Q1[2]} ,R2[11] ) ;
    _4R2Q_R4 _4R2Q_R4_13( {R1[13],R1[9],R1[5],R1[1] }, {Q1[8],Q1[4]} ,R2[13] ) ;
    _4R2Q_R4 _4R2Q_R4_15( {R1[15],R1[11],R1[7],R1[3] }, {Q1[10],Q1[6]} ,R2[15] ) ;
    _4R2Q_R4 _4R2Q_R4_17( {R1[17],R1[13],R1[9],R1[5] }, {Q1[12],Q1[8]} ,R2[17] ) ;
    _4R2Q_R4 _4R2Q_R4_19( {R1[19],R1[15],R1[11],R1[7] }, {Q1[14],Q1[10]} ,R2[19] ) ;
    _4R2Q_R4 _4R2Q_R4_21( {R1[21],R1[17],R1[13],R1[9] }, {Q1[16],Q1[12]} ,R2[21] ) ;
    _4R2Q_R4 _4R2Q_R4_23( {R1[23],R1[19],R1[15],R1[11] }, {Q1[18],Q1[14]} ,R2[23] ) ;
    _4R2Q_R4 _4R2Q_R4_25( {R1[25],R1[21],R1[17],R1[13] }, {Q1[20],Q1[16]} ,R2[25] ) ;
    _4R2Q_R4 _4R2Q_R4_27( {R1[27],R1[23],R1[19],R1[15] }, {Q1[22],Q1[18]} ,R2[27] ) ;
    _4R2Q_R4 _4R2Q_R4_29( {R1[29],R1[25],R1[21],R1[17] }, {Q1[24],Q1[20]} ,R2[29] ) ;
    _4R2Q_R4 _4R2Q_R4_31( {R1[31],R1[27],R1[23],R1[19] }, {Q1[26],Q1[22]} ,R2[31] ) ;
    _4R2Q_R4 _4R2Q_R4_33( {R1[33],R1[29],R1[25],R1[21] }, {Q1[28],Q1[24]} ,R2[33] ) ;
    _4R2Q_R4 _4R2Q_R4_35( {R1[35],R1[31],R1[27],R1[23] }, {Q1[30],Q1[26]} ,R2[35] ) ;
    _4R2Q_R4 _4R2Q_R4_37( {R1[37],R1[33],R1[29],R1[25] }, {Q1[32],Q1[28]} ,R2[37] ) ;
    _4R2Q_R4 _4R2Q_R4_39( {R1[39],R1[35],R1[31],R1[27] }, {Q1[34],Q1[30]} ,R2[39] ) ;
    _4R2Q_R4 _4R2Q_R4_41( {R1[41],R1[37],R1[33],R1[29] }, {Q1[36],Q1[32]} ,R2[41] ) ;
    _4R2Q_R4 _4R2Q_R4_43( {R1[43],R1[39],R1[35],R1[31] }, {Q1[38],Q1[34]} ,R2[43] ) ;
    _4R2Q_R4 _4R2Q_R4_45( {R1[45],R1[41],R1[37],R1[33] }, {Q1[40],Q1[36]} ,R2[45] ) ;
    _4R2Q_R4 _4R2Q_R4_47( {R1[47],R1[43],R1[39],R1[35] }, {Q1[42],Q1[38]} ,R2[47] ) ;
    _4R2Q_R4 _4R2Q_R4_49( {R1[49],R1[45],R1[41],R1[37] }, {Q1[44],Q1[40]} ,R2[49] ) ;
    _4R2Q_R4 _4R2Q_R4_51( {R1[51],R1[47],R1[43],R1[39] }, {Q1[46],Q1[42]} ,R2[51] ) ;
    _4R2Q_R4 _4R2Q_R4_53( {R1[53],R1[49],R1[45],R1[41] }, {Q1[48],Q1[44]} ,R2[53] ) ;
    _4R2Q_R4 _4R2Q_R4_55( {R1[55],R1[51],R1[47],R1[43] }, {Q1[50],Q1[46]} ,R2[55] ) ;
    _4R2Q_R4 _4R2Q_R4_57( {R1[57],R1[53],R1[49],R1[45] }, {Q1[52],Q1[48]} ,R2[57] ) ;
    _4R2Q_R4 _4R2Q_R4_59( {R1[59],R1[55],R1[51],R1[47] }, {Q1[54],Q1[50]} ,R2[59] ) ;
    _4R2Q_R4 _4R2Q_R4_61( {R1[61],R1[57],R1[53],R1[49] }, {Q1[56],Q1[52]} ,R2[61] ) ;
    _4R2Q_R4 _4R2Q_R4_63( {R1[63],R1[59],R1[55],R1[51] }, {Q1[58],Q1[54]} ,R2[63] ) ;

    _1R4Q_Q4 _1R4Q_Q4_0(R1[53], {Q1[0],Q1[60],Q1[56],Q1[52]}, Q2[0] ) ;
    _1R4Q_Q4 _1R4Q_Q4_2(R1[55], {Q1[2],Q1[62],Q1[58],Q1[54]}, Q2[2] ) ;
    _1R4Q_Q4 _1R4Q_Q4_4(R1[57], {Q1[4],Q1[0],Q1[60],Q1[56]}, Q2[4] ) ;
    _1R4Q_Q4 _1R4Q_Q4_6(R1[59], {Q1[6],Q1[2],Q1[62],Q1[58]}, Q2[6] ) ;
    _1R4Q_Q4 _1R4Q_Q4_8(R1[61], {Q1[8],Q1[4],Q1[0],Q1[60]}, Q2[8] ) ;
    _1R4Q_Q4 _1R4Q_Q4_10(R1[63], {Q1[10],Q1[6],Q1[2],Q1[62]}, Q2[10] ) ;
    _1R4Q_Q4 _1R4Q_Q4_12(R1[1], {Q1[12],Q1[8],Q1[4],Q1[0]}, Q2[12] ) ;
    _1R4Q_Q4 _1R4Q_Q4_14(R1[3], {Q1[14],Q1[10],Q1[6],Q1[2]}, Q2[14] ) ;
    _1R4Q_Q4 _1R4Q_Q4_16(R1[5], {Q1[16],Q1[12],Q1[8],Q1[4]}, Q2[16] ) ;
    _1R4Q_Q4 _1R4Q_Q4_18(R1[7], {Q1[18],Q1[14],Q1[10],Q1[6]}, Q2[18] ) ;
    _1R4Q_Q4 _1R4Q_Q4_20(R1[9], {Q1[20],Q1[16],Q1[12],Q1[8]}, Q2[20] ) ;
    _1R4Q_Q4 _1R4Q_Q4_22(R1[11], {Q1[22],Q1[18],Q1[14],Q1[10]}, Q2[22] ) ;
    _1R4Q_Q4 _1R4Q_Q4_24(R1[13], {Q1[24],Q1[20],Q1[16],Q1[12]}, Q2[24] ) ;
    _1R4Q_Q4 _1R4Q_Q4_26(R1[15], {Q1[26],Q1[22],Q1[18],Q1[14]}, Q2[26] ) ;
    _1R4Q_Q4 _1R4Q_Q4_28(R1[17], {Q1[28],Q1[24],Q1[20],Q1[16]}, Q2[28] ) ;
    _1R4Q_Q4 _1R4Q_Q4_30(R1[19], {Q1[30],Q1[26],Q1[22],Q1[18]}, Q2[30] ) ;
    _1R4Q_Q4 _1R4Q_Q4_32(R1[21], {Q1[32],Q1[28],Q1[24],Q1[20]}, Q2[32] ) ;
    _1R4Q_Q4 _1R4Q_Q4_34(R1[23], {Q1[34],Q1[30],Q1[26],Q1[22]}, Q2[34] ) ;
    _1R4Q_Q4 _1R4Q_Q4_36(R1[25], {Q1[36],Q1[32],Q1[28],Q1[24]}, Q2[36] ) ;
    _1R4Q_Q4 _1R4Q_Q4_38(R1[27], {Q1[38],Q1[34],Q1[30],Q1[26]}, Q2[38] ) ;
    _1R4Q_Q4 _1R4Q_Q4_40(R1[29], {Q1[40],Q1[36],Q1[32],Q1[28]}, Q2[40] ) ;
    _1R4Q_Q4 _1R4Q_Q4_42(R1[31], {Q1[42],Q1[38],Q1[34],Q1[30]}, Q2[42] ) ;
    _1R4Q_Q4 _1R4Q_Q4_44(R1[33], {Q1[44],Q1[40],Q1[36],Q1[32]}, Q2[44] ) ;
    _1R4Q_Q4 _1R4Q_Q4_46(R1[35], {Q1[46],Q1[42],Q1[38],Q1[34]}, Q2[46] ) ;
    _1R4Q_Q4 _1R4Q_Q4_48(R1[37], {Q1[48],Q1[44],Q1[40],Q1[36]}, Q2[48] ) ;
    _1R4Q_Q4 _1R4Q_Q4_50(R1[39], {Q1[50],Q1[46],Q1[42],Q1[38]}, Q2[50] ) ;
    _1R4Q_Q4 _1R4Q_Q4_52(R1[41], {Q1[52],Q1[48],Q1[44],Q1[40]}, Q2[52] ) ;
    _1R4Q_Q4 _1R4Q_Q4_54(R1[43], {Q1[54],Q1[50],Q1[46],Q1[42]}, Q2[54] ) ;
    _1R4Q_Q4 _1R4Q_Q4_56(R1[45], {Q1[56],Q1[52],Q1[48],Q1[44]}, Q2[56] ) ;
    _1R4Q_Q4 _1R4Q_Q4_58(R1[47], {Q1[58],Q1[54],Q1[50],Q1[46]}, Q2[58] ) ;
    _1R4Q_Q4 _1R4Q_Q4_60(R1[49], {Q1[60],Q1[56],Q1[52],Q1[48]}, Q2[60] ) ;
    _1R4Q_Q4 _1R4Q_Q4_62(R1[51], {Q1[62],Q1[58],Q1[54],Q1[50]}, Q2[62] ) ;

    _4R2Q_R4 _4R2Q_R4_65( {R2[1],R2[49],R2[33],R2[17] }, {Q2[44],Q2[28]} ,R3[1] ) ;
    _4R2Q_R4 _4R2Q_R4_67( {R2[3],R2[51],R2[35],R2[19] }, {Q2[46],Q2[30]} ,R3[3] ) ;
    _4R2Q_R4 _4R2Q_R4_69( {R2[5],R2[53],R2[37],R2[21] }, {Q2[48],Q2[32]} ,R3[5] ) ;
    _4R2Q_R4 _4R2Q_R4_71( {R2[7],R2[55],R2[39],R2[23] }, {Q2[50],Q2[34]} ,R3[7] ) ;
    _4R2Q_R4 _4R2Q_R4_73( {R2[9],R2[57],R2[41],R2[25] }, {Q2[52],Q2[36]} ,R3[9] ) ;
    _4R2Q_R4 _4R2Q_R4_75( {R2[11],R2[59],R2[43],R2[27] }, {Q2[54],Q2[38]} ,R3[11] ) ;
    _4R2Q_R4 _4R2Q_R4_77( {R2[13],R2[61],R2[45],R2[29] }, {Q2[56],Q2[40]} ,R3[13] ) ;
    _4R2Q_R4 _4R2Q_R4_79( {R2[15],R2[63],R2[47],R2[31] }, {Q2[58],Q2[42]} ,R3[15] ) ;
    _4R2Q_R4 _4R2Q_R4_81( {R2[17],R2[1],R2[49],R2[33] }, {Q2[60],Q2[44]} ,R3[17] ) ;
    _4R2Q_R4 _4R2Q_R4_83( {R2[19],R2[3],R2[51],R2[35] }, {Q2[62],Q2[46]} ,R3[19] ) ;
    _4R2Q_R4 _4R2Q_R4_85( {R2[21],R2[5],R2[53],R2[37] }, {Q2[0],Q2[48]} ,R3[21] ) ;
    _4R2Q_R4 _4R2Q_R4_87( {R2[23],R2[7],R2[55],R2[39] }, {Q2[2],Q2[50]} ,R3[23] ) ;
    _4R2Q_R4 _4R2Q_R4_89( {R2[25],R2[9],R2[57],R2[41] }, {Q2[4],Q2[52]} ,R3[25] ) ;
    _4R2Q_R4 _4R2Q_R4_91( {R2[27],R2[11],R2[59],R2[43] }, {Q2[6],Q2[54]} ,R3[27] ) ;
    _4R2Q_R4 _4R2Q_R4_93( {R2[29],R2[13],R2[61],R2[45] }, {Q2[8],Q2[56]} ,R3[29] ) ;
    _4R2Q_R4 _4R2Q_R4_95( {R2[31],R2[15],R2[63],R2[47] }, {Q2[10],Q2[58]} ,R3[31] ) ;
    _4R2Q_R4 _4R2Q_R4_97( {R2[33],R2[17],R2[1],R2[49] }, {Q2[12],Q2[60]} ,R3[33] ) ;
    _4R2Q_R4 _4R2Q_R4_99( {R2[35],R2[19],R2[3],R2[51] }, {Q2[14],Q2[62]} ,R3[35] ) ;
    _4R2Q_R4 _4R2Q_R4_101( {R2[37],R2[21],R2[5],R2[53] }, {Q2[16],Q2[0]} ,R3[37] ) ;
    _4R2Q_R4 _4R2Q_R4_103( {R2[39],R2[23],R2[7],R2[55] }, {Q2[18],Q2[2]} ,R3[39] ) ;
    _4R2Q_R4 _4R2Q_R4_105( {R2[41],R2[25],R2[9],R2[57] }, {Q2[20],Q2[4]} ,R3[41] ) ;
    _4R2Q_R4 _4R2Q_R4_107( {R2[43],R2[27],R2[11],R2[59] }, {Q2[22],Q2[6]} ,R3[43] ) ;
    _4R2Q_R4 _4R2Q_R4_109( {R2[45],R2[29],R2[13],R2[61] }, {Q2[24],Q2[8]} ,R3[45] ) ;
    _4R2Q_R4 _4R2Q_R4_111( {R2[47],R2[31],R2[15],R2[63] }, {Q2[26],Q2[10]} ,R3[47] ) ;
    _4R2Q_R4 _4R2Q_R4_113( {R2[49],R2[33],R2[17],R2[1] }, {Q2[28],Q2[12]} ,R3[49] ) ;
    _4R2Q_R4 _4R2Q_R4_115( {R2[51],R2[35],R2[19],R2[3] }, {Q2[30],Q2[14]} ,R3[51] ) ;
    _4R2Q_R4 _4R2Q_R4_117( {R2[53],R2[37],R2[21],R2[5] }, {Q2[32],Q2[16]} ,R3[53] ) ;
    _4R2Q_R4 _4R2Q_R4_119( {R2[55],R2[39],R2[23],R2[7] }, {Q2[34],Q2[18]} ,R3[55] ) ;
    _4R2Q_R4 _4R2Q_R4_121( {R2[57],R2[41],R2[25],R2[9] }, {Q2[36],Q2[20]} ,R3[57] ) ;
    _4R2Q_R4 _4R2Q_R4_123( {R2[59],R2[43],R2[27],R2[11] }, {Q2[38],Q2[22]} ,R3[59] ) ;
    _4R2Q_R4 _4R2Q_R4_125( {R2[61],R2[45],R2[29],R2[13] }, {Q2[40],Q2[24]} ,R3[61] ) ;
    _4R2Q_R4 _4R2Q_R4_127( {R2[63],R2[47],R2[31],R2[15] }, {Q2[42],Q2[26]} ,R3[63] ) ;

    _D64_1 _D64_1_1( {p[1],p[0],p[63]}, {g[1],g[0]}, D1[1] ) ;
    _D64_1 _D64_1_3( {p[3],p[2],p[1]}, {g[3],g[2]}, D1[3] ) ;
    _D64_1 _D64_1_5( {p[5],p[4],p[3]}, {g[5],g[4]}, D1[5] ) ;
    _D64_1 _D64_1_7( {p[7],p[6],p[5]}, {g[7],g[6]}, D1[7] ) ;
    _D64_1 _D64_1_9( {p[9],p[8],p[7]}, {g[9],g[8]}, D1[9] ) ;
    _D64_1 _D64_1_11( {p[11],p[10],p[9]}, {g[11],g[10]}, D1[11] ) ;
    _D64_1 _D64_1_13( {p[13],p[12],p[11]}, {g[13],g[12]}, D1[13] ) ;
    _D64_1 _D64_1_15( {p[15],p[14],p[13]}, {g[15],g[14]}, D1[15] ) ;
    _D64_1 _D64_1_17( {p[17],p[16],p[15]}, {g[17],g[16]}, D1[17] ) ;
    _D64_1 _D64_1_19( {p[19],p[18],p[17]}, {g[19],g[18]}, D1[19] ) ;
    _D64_1 _D64_1_21( {p[21],p[20],p[19]}, {g[21],g[20]}, D1[21] ) ;
    _D64_1 _D64_1_23( {p[23],p[22],p[21]}, {g[23],g[22]}, D1[23] ) ;
    _D64_1 _D64_1_25( {p[25],p[24],p[23]}, {g[25],g[24]}, D1[25] ) ;
    _D64_1 _D64_1_27( {p[27],p[26],p[25]}, {g[27],g[26]}, D1[27] ) ;
    _D64_1 _D64_1_29( {p[29],p[28],p[27]}, {g[29],g[28]}, D1[29] ) ;
    _D64_1 _D64_1_31( {p[31],p[30],p[29]}, {g[31],g[30]}, D1[31] ) ;
    _D64_1 _D64_1_33( {p[33],p[32],p[31]}, {g[33],g[32]}, D1[33] ) ;
    _D64_1 _D64_1_35( {p[35],p[34],p[33]}, {g[35],g[34]}, D1[35] ) ;
    _D64_1 _D64_1_37( {p[37],p[36],p[35]}, {g[37],g[36]}, D1[37] ) ;
    _D64_1 _D64_1_39( {p[39],p[38],p[37]}, {g[39],g[38]}, D1[39] ) ;
    _D64_1 _D64_1_41( {p[41],p[40],p[39]}, {g[41],g[40]}, D1[41] ) ;
    _D64_1 _D64_1_43( {p[43],p[42],p[41]}, {g[43],g[42]}, D1[43] ) ;
    _D64_1 _D64_1_45( {p[45],p[44],p[43]}, {g[45],g[44]}, D1[45] ) ;
    _D64_1 _D64_1_47( {p[47],p[46],p[45]}, {g[47],g[46]}, D1[47] ) ;
    _D64_1 _D64_1_49( {p[49],p[48],p[47]}, {g[49],g[48]}, D1[49] ) ;
    _D64_1 _D64_1_51( {p[51],p[50],p[49]}, {g[51],g[50]}, D1[51] ) ;
    _D64_1 _D64_1_53( {p[53],p[52],p[51]}, {g[53],g[52]}, D1[53] ) ;
    _D64_1 _D64_1_55( {p[55],p[54],p[53]}, {g[55],g[54]}, D1[55] ) ;
    _D64_1 _D64_1_57( {p[57],p[56],p[55]}, {g[57],g[56]}, D1[57] ) ;
    _D64_1 _D64_1_59( {p[59],p[58],p[57]}, {g[59],g[58]}, D1[59] ) ;
    _D64_1 _D64_1_61( {p[61],p[60],p[59]}, {g[61],g[60]}, D1[61] ) ;
    _D64_1 _D64_1_63( {p[63],p[62],p[61]}, {g[63],g[62]}, D1[63] ) ;

    _D64_2 _D64_2_1(D1[1] ,R1[1] ,Q1[0] ,D2[1] ) ;
    _D64_2 _D64_2_3(D1[3] ,R1[3] ,Q1[2] ,D2[3] ) ;
    _D64_2 _D64_2_5(D1[5] ,R1[5] ,Q1[4] ,D2[5] ) ;
    _D64_2 _D64_2_7(D1[7] ,R1[7] ,Q1[6] ,D2[7] ) ;
    _D64_2 _D64_2_9(D1[9] ,R1[9] ,Q1[8] ,D2[9] ) ;
    _D64_2 _D64_2_11(D1[11] ,R1[11] ,Q1[10] ,D2[11] ) ;
    _D64_2 _D64_2_13(D1[13] ,R1[13] ,Q1[12] ,D2[13] ) ;
    _D64_2 _D64_2_15(D1[15] ,R1[15] ,Q1[14] ,D2[15] ) ;
    _D64_2 _D64_2_17(D1[17] ,R1[17] ,Q1[16] ,D2[17] ) ;
    _D64_2 _D64_2_19(D1[19] ,R1[19] ,Q1[18] ,D2[19] ) ;
    _D64_2 _D64_2_21(D1[21] ,R1[21] ,Q1[20] ,D2[21] ) ;
    _D64_2 _D64_2_23(D1[23] ,R1[23] ,Q1[22] ,D2[23] ) ;
    _D64_2 _D64_2_25(D1[25] ,R1[25] ,Q1[24] ,D2[25] ) ;
    _D64_2 _D64_2_27(D1[27] ,R1[27] ,Q1[26] ,D2[27] ) ;
    _D64_2 _D64_2_29(D1[29] ,R1[29] ,Q1[28] ,D2[29] ) ;
    _D64_2 _D64_2_31(D1[31] ,R1[31] ,Q1[30] ,D2[31] ) ;
    _D64_2 _D64_2_33(D1[33] ,R1[33] ,Q1[32] ,D2[33] ) ;
    _D64_2 _D64_2_35(D1[35] ,R1[35] ,Q1[34] ,D2[35] ) ;
    _D64_2 _D64_2_37(D1[37] ,R1[37] ,Q1[36] ,D2[37] ) ;
    _D64_2 _D64_2_39(D1[39] ,R1[39] ,Q1[38] ,D2[39] ) ;
    _D64_2 _D64_2_41(D1[41] ,R1[41] ,Q1[40] ,D2[41] ) ;
    _D64_2 _D64_2_43(D1[43] ,R1[43] ,Q1[42] ,D2[43] ) ;
    _D64_2 _D64_2_45(D1[45] ,R1[45] ,Q1[44] ,D2[45] ) ;
    _D64_2 _D64_2_47(D1[47] ,R1[47] ,Q1[46] ,D2[47] ) ;
    _D64_2 _D64_2_49(D1[49] ,R1[49] ,Q1[48] ,D2[49] ) ;
    _D64_2 _D64_2_51(D1[51] ,R1[51] ,Q1[50] ,D2[51] ) ;
    _D64_2 _D64_2_53(D1[53] ,R1[53] ,Q1[52] ,D2[53] ) ;
    _D64_2 _D64_2_55(D1[55] ,R1[55] ,Q1[54] ,D2[55] ) ;
    _D64_2 _D64_2_57(D1[57] ,R1[57] ,Q1[56] ,D2[57] ) ;
    _D64_2 _D64_2_59(D1[59] ,R1[59] ,Q1[58] ,D2[59] ) ;
    _D64_2 _D64_2_61(D1[61] ,R1[61] ,Q1[60] ,D2[61] ) ;
    _D64_2 _D64_2_63(D1[63] ,R1[63] ,Q1[62] ,D2[63] ) ;

    _D64_2 _D64_2_65(D2[1] ,R2[1] ,Q2[60] ,D3[1] ) ;
    _D64_2 _D64_2_67(D2[3] ,R2[3] ,Q2[62] ,D3[3] ) ;
    _D64_2 _D64_2_69(D2[5] ,R2[5] ,Q2[0] ,D3[5] ) ;
    _D64_2 _D64_2_71(D2[7] ,R2[7] ,Q2[2] ,D3[7] ) ;
    _D64_2 _D64_2_73(D2[9] ,R2[9] ,Q2[4] ,D3[9] ) ;
    _D64_2 _D64_2_75(D2[11] ,R2[11] ,Q2[6] ,D3[11] ) ;
    _D64_2 _D64_2_77(D2[13] ,R2[13] ,Q2[8] ,D3[13] ) ;
    _D64_2 _D64_2_79(D2[15] ,R2[15] ,Q2[10] ,D3[15] ) ;
    _D64_2 _D64_2_81(D2[17] ,R2[17] ,Q2[12] ,D3[17] ) ;
    _D64_2 _D64_2_83(D2[19] ,R2[19] ,Q2[14] ,D3[19] ) ;
    _D64_2 _D64_2_85(D2[21] ,R2[21] ,Q2[16] ,D3[21] ) ;
    _D64_2 _D64_2_87(D2[23] ,R2[23] ,Q2[18] ,D3[23] ) ;
    _D64_2 _D64_2_89(D2[25] ,R2[25] ,Q2[20] ,D3[25] ) ;
    _D64_2 _D64_2_91(D2[27] ,R2[27] ,Q2[22] ,D3[27] ) ;
    _D64_2 _D64_2_93(D2[29] ,R2[29] ,Q2[24] ,D3[29] ) ;
    _D64_2 _D64_2_95(D2[31] ,R2[31] ,Q2[26] ,D3[31] ) ;
    _D64_2 _D64_2_97(D2[33] ,R2[33] ,Q2[28] ,D3[33] ) ;
    _D64_2 _D64_2_99(D2[35] ,R2[35] ,Q2[30] ,D3[35] ) ;
    _D64_2 _D64_2_101(D2[37] ,R2[37] ,Q2[32] ,D3[37] ) ;
    _D64_2 _D64_2_103(D2[39] ,R2[39] ,Q2[34] ,D3[39] ) ;
    _D64_2 _D64_2_105(D2[41] ,R2[41] ,Q2[36] ,D3[41] ) ;
    _D64_2 _D64_2_107(D2[43] ,R2[43] ,Q2[38] ,D3[43] ) ;
    _D64_2 _D64_2_109(D2[45] ,R2[45] ,Q2[40] ,D3[45] ) ;
    _D64_2 _D64_2_111(D2[47] ,R2[47] ,Q2[42] ,D3[47] ) ;
    _D64_2 _D64_2_113(D2[49] ,R2[49] ,Q2[44] ,D3[49] ) ;
    _D64_2 _D64_2_115(D2[51] ,R2[51] ,Q2[46] ,D3[51] ) ;
    _D64_2 _D64_2_117(D2[53] ,R2[53] ,Q2[48] ,D3[53] ) ;
    _D64_2 _D64_2_119(D2[55] ,R2[55] ,Q2[50] ,D3[55] ) ;
    _D64_2 _D64_2_121(D2[57] ,R2[57] ,Q2[52] ,D3[57] ) ;
    _D64_2 _D64_2_123(D2[59] ,R2[59] ,Q2[54] ,D3[59] ) ;
    _D64_2 _D64_2_125(D2[61] ,R2[61] ,Q2[56] ,D3[61] ) ;
    _D64_2 _D64_2_127(D2[63] ,R2[63] ,Q2[58] ,D3[63] ) ;

    _Jsum_sparse2 _Jsum_sparse2_0( g[0] , p[0] , R3[63], D3[63] , {x[1],x[0]} , {sum[1],sum[0]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_2( g[2] , p[2] , R3[1], D3[1] , {x[3],x[2]} , {sum[3],sum[2]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_4( g[4] , p[4] , R3[3], D3[3] , {x[5],x[4]} , {sum[5],sum[4]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_6( g[6] , p[6] , R3[5], D3[5] , {x[7],x[6]} , {sum[7],sum[6]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_8( g[8] , p[8] , R3[7], D3[7] , {x[9],x[8]} , {sum[9],sum[8]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_10( g[10] , p[10] , R3[9], D3[9] , {x[11],x[10]} , {sum[11],sum[10]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_12( g[12] , p[12] , R3[11], D3[11] , {x[13],x[12]} , {sum[13],sum[12]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_14( g[14] , p[14] , R3[13], D3[13] , {x[15],x[14]} , {sum[15],sum[14]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_16( g[16] , p[16] , R3[15], D3[15] , {x[17],x[16]} , {sum[17],sum[16]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_18( g[18] , p[18] , R3[17], D3[17] , {x[19],x[18]} , {sum[19],sum[18]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_20( g[20] , p[20] , R3[19], D3[19] , {x[21],x[20]} , {sum[21],sum[20]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_22( g[22] , p[22] , R3[21], D3[21] , {x[23],x[22]} , {sum[23],sum[22]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_24( g[24] , p[24] , R3[23], D3[23] , {x[25],x[24]} , {sum[25],sum[24]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_26( g[26] , p[26] , R3[25], D3[25] , {x[27],x[26]} , {sum[27],sum[26]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_28( g[28] , p[28] , R3[27], D3[27] , {x[29],x[28]} , {sum[29],sum[28]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_30( g[30] , p[30] , R3[29], D3[29] , {x[31],x[30]} , {sum[31],sum[30]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_32( g[32] , p[32] , R3[31], D3[31] , {x[33],x[32]} , {sum[33],sum[32]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_34( g[34] , p[34] , R3[33], D3[33] , {x[35],x[34]} , {sum[35],sum[34]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_36( g[36] , p[36] , R3[35], D3[35] , {x[37],x[36]} , {sum[37],sum[36]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_38( g[38] , p[38] , R3[37], D3[37] , {x[39],x[38]} , {sum[39],sum[38]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_40( g[40] , p[40] , R3[39], D3[39] , {x[41],x[40]} , {sum[41],sum[40]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_42( g[42] , p[42] , R3[41], D3[41] , {x[43],x[42]} , {sum[43],sum[42]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_44( g[44] , p[44] , R3[43], D3[43] , {x[45],x[44]} , {sum[45],sum[44]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_46( g[46] , p[46] , R3[45], D3[45] , {x[47],x[46]} , {sum[47],sum[46]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_48( g[48] , p[48] , R3[47], D3[47] , {x[49],x[48]} , {sum[49],sum[48]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_50( g[50] , p[50] , R3[49], D3[49] , {x[51],x[50]} , {sum[51],sum[50]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_52( g[52] , p[52] , R3[51], D3[51] , {x[53],x[52]} , {sum[53],sum[52]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_54( g[54] , p[54] , R3[53], D3[53] , {x[55],x[54]} , {sum[55],sum[54]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_56( g[56] , p[56] , R3[55], D3[55] , {x[57],x[56]} , {sum[57],sum[56]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_58( g[58] , p[58] , R3[57], D3[57] , {x[59],x[58]} , {sum[59],sum[58]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_60( g[60] , p[60] , R3[59], D3[59] , {x[61],x[60]} , {sum[61],sum[60]} ) ;
    _Jsum_sparse2 _Jsum_sparse2_62( g[62] , p[62] , R3[61], D3[61] , {x[63],x[62]} , {sum[63],sum[62]} ) ;

endmodule
